magic
tech sky130A
magscale 1 2
timestamp 1614532229
<< obsli1 >>
rect 1104 2159 21712 22321
<< obsm1 >>
rect 566 2128 22158 22352
<< metal2 >>
rect 2042 24202 2098 25002
rect 4802 24202 4858 25002
rect 7746 24202 7802 25002
rect 10690 24202 10746 25002
rect 13450 24202 13506 25002
rect 16394 24202 16450 25002
rect 19338 24202 19394 25002
rect 22098 24202 22154 25002
rect 570 0 626 800
rect 3330 0 3386 800
rect 6274 0 6330 800
rect 9218 0 9274 800
rect 11978 0 12034 800
rect 14922 0 14978 800
rect 17866 0 17922 800
rect 20626 0 20682 800
<< obsm2 >>
rect 572 24146 1986 24202
rect 2154 24146 4746 24202
rect 4914 24146 7690 24202
rect 7858 24146 10634 24202
rect 10802 24146 13394 24202
rect 13562 24146 16338 24202
rect 16506 24146 19282 24202
rect 19450 24146 22042 24202
rect 572 856 22152 24146
rect 682 800 3274 856
rect 3442 800 6218 856
rect 6386 800 9162 856
rect 9330 800 11922 856
rect 12090 800 14866 856
rect 15034 800 17810 856
rect 17978 800 20570 856
rect 20738 800 22152 856
<< metal3 >>
rect 0 22040 800 22160
rect 22058 19864 22858 19984
rect 0 17688 800 17808
rect 22058 15512 22858 15632
rect 0 13608 800 13728
rect 22058 11160 22858 11280
rect 0 9256 800 9376
rect 22058 7080 22858 7200
rect 0 4904 800 5024
rect 22058 2728 22858 2848
<< obsm3 >>
rect 800 22240 22058 22337
rect 880 21960 22058 22240
rect 800 20064 22058 21960
rect 800 19784 21978 20064
rect 800 17888 22058 19784
rect 880 17608 22058 17888
rect 800 15712 22058 17608
rect 800 15432 21978 15712
rect 800 13808 22058 15432
rect 880 13528 22058 13808
rect 800 11360 22058 13528
rect 800 11080 21978 11360
rect 800 9456 22058 11080
rect 880 9176 22058 9456
rect 800 7280 22058 9176
rect 800 7000 21978 7280
rect 800 5104 22058 7000
rect 880 4824 22058 5104
rect 800 2928 22058 4824
rect 800 2648 21978 2928
rect 800 2143 22058 2648
<< metal4 >>
rect 4379 2128 4699 22352
rect 7813 2128 8133 22352
rect 11248 2128 11568 22352
rect 14683 2128 15003 22352
rect 18117 2128 18437 22352
<< obsm4 >>
rect 4779 2128 7733 22352
rect 8213 2128 11168 22352
rect 11648 2128 14603 22352
<< metal5 >>
rect 1104 18741 21712 19061
rect 1104 15387 21712 15707
rect 1104 12032 21712 12352
rect 1104 8677 21712 8997
rect 1104 5323 21712 5643
<< obsm5 >>
rect 1104 12672 21712 15067
rect 1104 9317 21712 11712
rect 1104 5963 21712 8357
<< labels >>
rlabel metal2 s 2042 24202 2098 25002 6 ci
port 1 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 co
port 2 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 i0[0]
port 3 nsew signal input
rlabel metal2 s 570 0 626 800 6 i0[1]
port 4 nsew signal input
rlabel metal2 s 7746 24202 7802 25002 6 i0[2]
port 5 nsew signal input
rlabel metal3 s 22058 7080 22858 7200 6 i0[3]
port 6 nsew signal input
rlabel metal3 s 22058 15512 22858 15632 6 i0[4]
port 7 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 i0[5]
port 8 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 i0[6]
port 9 nsew signal input
rlabel metal2 s 19338 24202 19394 25002 6 i0[7]
port 10 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 i1[0]
port 11 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 i1[1]
port 12 nsew signal input
rlabel metal3 s 22058 19864 22858 19984 6 i1[2]
port 13 nsew signal input
rlabel metal3 s 22058 11160 22858 11280 6 i1[3]
port 14 nsew signal input
rlabel metal2 s 22098 24202 22154 25002 6 i1[4]
port 15 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 i1[5]
port 16 nsew signal input
rlabel metal2 s 10690 24202 10746 25002 6 i1[6]
port 17 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 i1[7]
port 18 nsew signal input
rlabel metal2 s 4802 24202 4858 25002 6 s[0]
port 19 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 s[1]
port 20 nsew signal output
rlabel metal2 s 13450 24202 13506 25002 6 s[2]
port 21 nsew signal output
rlabel metal3 s 22058 2728 22858 2848 6 s[3]
port 22 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 s[4]
port 23 nsew signal output
rlabel metal2 s 16394 24202 16450 25002 6 s[5]
port 24 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 s[6]
port 25 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 s[7]
port 26 nsew signal output
rlabel metal4 s 18117 2128 18437 22352 6 VPWR
port 27 nsew power bidirectional
rlabel metal4 s 11248 2128 11568 22352 6 VPWR
port 28 nsew power bidirectional
rlabel metal4 s 4379 2128 4699 22352 6 VPWR
port 29 nsew power bidirectional
rlabel metal5 s 1104 18741 21712 19061 6 VPWR
port 30 nsew power bidirectional
rlabel metal5 s 1104 12032 21712 12352 6 VPWR
port 31 nsew power bidirectional
rlabel metal5 s 1104 5323 21712 5643 6 VPWR
port 32 nsew power bidirectional
rlabel metal4 s 14683 2128 15003 22352 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 7813 2128 8133 22352 6 VGND
port 34 nsew ground bidirectional
rlabel metal5 s 1104 15387 21712 15707 6 VGND
port 35 nsew ground bidirectional
rlabel metal5 s 1104 8677 21712 8997 6 VGND
port 36 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22858 25002
string LEFview TRUE
<< end >>
