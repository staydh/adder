magic
tech sky130A
magscale 1 2
timestamp 1616762085
<< checkpaint >>
rect -3932 -3932 26790 28934
<< viali >>
rect 19349 21505 19383 21539
rect 19441 21437 19475 21471
rect 19993 21437 20027 21471
rect 20177 21437 20211 21471
rect 20453 21301 20487 21335
rect 19073 21097 19107 21131
rect 19441 20961 19475 20995
rect 19809 20961 19843 20995
rect 19993 20961 20027 20995
rect 19533 20893 19567 20927
rect 20361 20485 20395 20519
rect 19441 20349 19475 20383
rect 19533 20349 19567 20383
rect 19901 20349 19935 20383
rect 19993 20349 20027 20383
rect 19533 19873 19567 19907
rect 19441 19805 19475 19839
rect 19717 19669 19751 19703
rect 18889 19261 18923 19295
rect 19001 19261 19035 19295
rect 19441 19193 19475 19227
rect 18889 18921 18923 18955
rect 19257 18785 19291 18819
rect 19625 18785 19659 18819
rect 19349 18717 19383 18751
rect 19533 18717 19567 18751
rect 18797 18173 18831 18207
rect 18889 18173 18923 18207
rect 19257 18173 19291 18207
rect 19349 18173 19383 18207
rect 19809 18037 19843 18071
rect 19901 17765 19935 17799
rect 18613 17697 18647 17731
rect 18797 17697 18831 17731
rect 19349 17697 19383 17731
rect 19533 17697 19567 17731
rect 19441 17289 19475 17323
rect 19257 17085 19291 17119
rect 16405 16745 16439 16779
rect 16221 16609 16255 16643
rect 15761 16201 15795 16235
rect 16221 16065 16255 16099
rect 16405 16065 16439 16099
rect 16129 15997 16163 16031
rect 16497 15997 16531 16031
rect 19073 15657 19107 15691
rect 15761 15521 15795 15555
rect 16313 15521 16347 15555
rect 16497 15521 16531 15555
rect 17785 15521 17819 15555
rect 18889 15521 18923 15555
rect 15669 15453 15703 15487
rect 16773 15317 16807 15351
rect 17969 15317 18003 15351
rect 16129 15113 16163 15147
rect 15853 14909 15887 14943
rect 15945 14909 15979 14943
rect 17601 14501 17635 14535
rect 13369 14433 13403 14467
rect 16497 14433 16531 14467
rect 16957 14433 16991 14467
rect 17049 14433 17083 14467
rect 16405 14365 16439 14399
rect 13553 14229 13587 14263
rect 14565 14025 14599 14059
rect 13001 13821 13035 13855
rect 13093 13821 13127 13855
rect 14381 13821 14415 13855
rect 13553 13753 13587 13787
rect 12909 13481 12943 13515
rect 13277 13345 13311 13379
rect 13645 13345 13679 13379
rect 13737 13345 13771 13379
rect 13369 13277 13403 13311
rect 13645 12733 13679 12767
rect 13737 12733 13771 12767
rect 14105 12733 14139 12767
rect 14197 12733 14231 12767
rect 15669 12733 15703 12767
rect 14749 12665 14783 12699
rect 15853 12597 15887 12631
rect 14013 12325 14047 12359
rect 12909 12257 12943 12291
rect 13461 12257 13495 12291
rect 13645 12257 13679 12291
rect 12725 12189 12759 12223
rect 13553 11849 13587 11883
rect 10517 11645 10551 11679
rect 13369 11645 13403 11679
rect 10701 11509 10735 11543
rect 10701 11305 10735 11339
rect 13553 11305 13587 11339
rect 10517 11169 10551 11203
rect 11621 11169 11655 11203
rect 13369 11169 13403 11203
rect 11805 11033 11839 11067
rect 9229 10761 9263 10795
rect 9045 10557 9079 10591
rect 10149 10557 10183 10591
rect 10241 10557 10275 10591
rect 10701 10489 10735 10523
rect 13001 10217 13035 10251
rect 10793 10081 10827 10115
rect 10885 10081 10919 10115
rect 11253 10081 11287 10115
rect 11345 10081 11379 10115
rect 12817 10081 12851 10115
rect 11897 10013 11931 10047
rect 11069 9673 11103 9707
rect 9965 9537 9999 9571
rect 10057 9469 10091 9503
rect 10517 9469 10551 9503
rect 10609 9469 10643 9503
rect 10057 9129 10091 9163
rect 7665 8993 7699 9027
rect 10425 8993 10459 9027
rect 10793 8993 10827 9027
rect 10517 8925 10551 8959
rect 10701 8925 10735 8959
rect 7849 8789 7883 8823
rect 7849 8585 7883 8619
rect 10701 8585 10735 8619
rect 2421 8517 2455 8551
rect 8953 8517 8987 8551
rect 2237 8381 2271 8415
rect 7665 8381 7699 8415
rect 8769 8381 8803 8415
rect 10517 8381 10551 8415
rect 6377 8041 6411 8075
rect 2237 7905 2271 7939
rect 4813 7905 4847 7939
rect 6193 7905 6227 7939
rect 7389 7905 7423 7939
rect 7297 7837 7331 7871
rect 2421 7701 2455 7735
rect 4997 7701 5031 7735
rect 7573 7701 7607 7735
rect 10057 7497 10091 7531
rect 7757 7361 7791 7395
rect 2237 7293 2271 7327
rect 3341 7293 3375 7327
rect 4813 7293 4847 7327
rect 7849 7293 7883 7327
rect 8309 7293 8343 7327
rect 8401 7293 8435 7327
rect 9873 7293 9907 7327
rect 2421 7157 2455 7191
rect 3525 7157 3559 7191
rect 4997 7157 5031 7191
rect 8861 7157 8895 7191
rect 8217 6953 8251 6987
rect 2237 6817 2271 6851
rect 4813 6817 4847 6851
rect 5917 6817 5951 6851
rect 7205 6817 7239 6851
rect 7757 6817 7791 6851
rect 7941 6817 7975 6851
rect 7021 6749 7055 6783
rect 2421 6613 2455 6647
rect 4997 6613 5031 6647
rect 6101 6613 6135 6647
rect 7205 6409 7239 6443
rect 1777 6273 1811 6307
rect 4813 6273 4847 6307
rect 7481 6273 7515 6307
rect 7849 6273 7883 6307
rect 1869 6205 1903 6239
rect 4721 6205 4755 6239
rect 5043 6205 5077 6239
rect 5273 6205 5307 6239
rect 7573 6205 7607 6239
rect 7941 6205 7975 6239
rect 2329 6137 2363 6171
rect 4353 6069 4387 6103
rect 7849 5865 7883 5899
rect 2053 5729 2087 5763
rect 2421 5729 2455 5763
rect 2605 5729 2639 5763
rect 4813 5729 4847 5763
rect 4997 5729 5031 5763
rect 5457 5729 5491 5763
rect 5549 5729 5583 5763
rect 7665 5729 7699 5763
rect 1869 5661 1903 5695
rect 6009 5593 6043 5627
rect 1685 5525 1719 5559
rect 5365 5321 5399 5355
rect 2053 5185 2087 5219
rect 2145 5117 2179 5151
rect 2605 5117 2639 5151
rect 2697 5117 2731 5151
rect 4353 5117 4387 5151
rect 4445 5117 4479 5151
rect 4905 5117 4939 5151
rect 5089 5117 5123 5151
rect 6837 5117 6871 5151
rect 3249 5049 3283 5083
rect 7021 4981 7055 5015
rect 1501 4709 1535 4743
rect 4997 4709 5031 4743
rect 2329 4641 2363 4675
rect 2513 4641 2547 4675
rect 4537 4641 4571 4675
rect 5825 4641 5859 4675
rect 6929 4641 6963 4675
rect 2053 4573 2087 4607
rect 4445 4573 4479 4607
rect 6009 4437 6043 4471
rect 7113 4437 7147 4471
rect 2237 4029 2271 4063
rect 3341 4029 3375 4063
rect 4813 4029 4847 4063
rect 2421 3893 2455 3927
rect 3525 3893 3559 3927
rect 4997 3893 5031 3927
rect 2421 3689 2455 3723
rect 4997 3689 5031 3723
rect 2237 3553 2271 3587
rect 4813 3553 4847 3587
rect 2421 3145 2455 3179
rect 3433 3145 3467 3179
rect 2237 2941 2271 2975
rect 3341 2941 3375 2975
rect 2053 2601 2087 2635
rect 1961 2465 1995 2499
<< metal1 >>
rect 1104 22330 21712 22352
rect 1104 22278 7851 22330
rect 7903 22278 7915 22330
rect 7967 22278 7979 22330
rect 8031 22278 8043 22330
rect 8095 22278 14720 22330
rect 14772 22278 14784 22330
rect 14836 22278 14848 22330
rect 14900 22278 14912 22330
rect 14964 22278 21712 22330
rect 1104 22256 21712 22278
rect 1104 21786 21712 21808
rect 1104 21734 4416 21786
rect 4468 21734 4480 21786
rect 4532 21734 4544 21786
rect 4596 21734 4608 21786
rect 4660 21734 11286 21786
rect 11338 21734 11350 21786
rect 11402 21734 11414 21786
rect 11466 21734 11478 21786
rect 11530 21734 18155 21786
rect 18207 21734 18219 21786
rect 18271 21734 18283 21786
rect 18335 21734 18347 21786
rect 18399 21734 21712 21786
rect 1104 21712 21712 21734
rect 19242 21496 19248 21548
rect 19300 21536 19306 21548
rect 19337 21539 19395 21545
rect 19337 21536 19349 21539
rect 19300 21508 19349 21536
rect 19300 21496 19306 21508
rect 19337 21505 19349 21508
rect 19383 21536 19395 21539
rect 19383 21508 19564 21536
rect 19383 21505 19395 21508
rect 19337 21499 19395 21505
rect 19429 21471 19487 21477
rect 19429 21437 19441 21471
rect 19475 21437 19487 21471
rect 19536 21468 19564 21508
rect 19981 21471 20039 21477
rect 19981 21468 19993 21471
rect 19536 21440 19993 21468
rect 19429 21431 19487 21437
rect 19981 21437 19993 21440
rect 20027 21437 20039 21471
rect 20162 21468 20168 21480
rect 20123 21440 20168 21468
rect 19981 21431 20039 21437
rect 19444 21400 19472 21431
rect 20162 21428 20168 21440
rect 20220 21428 20226 21480
rect 20180 21400 20208 21428
rect 19444 21372 20208 21400
rect 20438 21332 20444 21344
rect 20399 21304 20444 21332
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 1104 21242 21712 21264
rect 1104 21190 7851 21242
rect 7903 21190 7915 21242
rect 7967 21190 7979 21242
rect 8031 21190 8043 21242
rect 8095 21190 14720 21242
rect 14772 21190 14784 21242
rect 14836 21190 14848 21242
rect 14900 21190 14912 21242
rect 14964 21190 21712 21242
rect 1104 21168 21712 21190
rect 19058 21128 19064 21140
rect 19019 21100 19064 21128
rect 19058 21088 19064 21100
rect 19116 21088 19122 21140
rect 19242 20952 19248 21004
rect 19300 20992 19306 21004
rect 19429 20995 19487 21001
rect 19429 20992 19441 20995
rect 19300 20964 19441 20992
rect 19300 20952 19306 20964
rect 19429 20961 19441 20964
rect 19475 20961 19487 20995
rect 19429 20955 19487 20961
rect 19610 20952 19616 21004
rect 19668 20992 19674 21004
rect 19797 20995 19855 21001
rect 19797 20992 19809 20995
rect 19668 20964 19809 20992
rect 19668 20952 19674 20964
rect 19797 20961 19809 20964
rect 19843 20961 19855 20995
rect 19797 20955 19855 20961
rect 19886 20952 19892 21004
rect 19944 20992 19950 21004
rect 19981 20995 20039 21001
rect 19981 20992 19993 20995
rect 19944 20964 19993 20992
rect 19944 20952 19950 20964
rect 19981 20961 19993 20964
rect 20027 20992 20039 20995
rect 21358 20992 21364 21004
rect 20027 20964 21364 20992
rect 20027 20961 20039 20964
rect 19981 20955 20039 20961
rect 21358 20952 21364 20964
rect 21416 20952 21422 21004
rect 19518 20924 19524 20936
rect 19479 20896 19524 20924
rect 19518 20884 19524 20896
rect 19576 20884 19582 20936
rect 1104 20698 21712 20720
rect 1104 20646 4416 20698
rect 4468 20646 4480 20698
rect 4532 20646 4544 20698
rect 4596 20646 4608 20698
rect 4660 20646 11286 20698
rect 11338 20646 11350 20698
rect 11402 20646 11414 20698
rect 11466 20646 11478 20698
rect 11530 20646 18155 20698
rect 18207 20646 18219 20698
rect 18271 20646 18283 20698
rect 18335 20646 18347 20698
rect 18399 20646 21712 20698
rect 1104 20624 21712 20646
rect 20162 20476 20168 20528
rect 20220 20516 20226 20528
rect 20349 20519 20407 20525
rect 20349 20516 20361 20519
rect 20220 20488 20361 20516
rect 20220 20476 20226 20488
rect 20349 20485 20361 20488
rect 20395 20485 20407 20519
rect 20349 20479 20407 20485
rect 19429 20383 19487 20389
rect 19429 20349 19441 20383
rect 19475 20349 19487 20383
rect 19429 20343 19487 20349
rect 19521 20383 19579 20389
rect 19521 20349 19533 20383
rect 19567 20380 19579 20383
rect 19886 20380 19892 20392
rect 19567 20352 19892 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 19444 20312 19472 20343
rect 19886 20340 19892 20352
rect 19944 20340 19950 20392
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20380 20039 20383
rect 20714 20380 20720 20392
rect 20027 20352 20720 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 19610 20312 19616 20324
rect 19444 20284 19616 20312
rect 19610 20272 19616 20284
rect 19668 20312 19674 20324
rect 19996 20312 20024 20343
rect 20714 20340 20720 20352
rect 20772 20340 20778 20392
rect 19668 20284 20024 20312
rect 19668 20272 19674 20284
rect 1104 20154 21712 20176
rect 1104 20102 7851 20154
rect 7903 20102 7915 20154
rect 7967 20102 7979 20154
rect 8031 20102 8043 20154
rect 8095 20102 14720 20154
rect 14772 20102 14784 20154
rect 14836 20102 14848 20154
rect 14900 20102 14912 20154
rect 14964 20102 21712 20154
rect 1104 20080 21712 20102
rect 19521 19907 19579 19913
rect 19521 19873 19533 19907
rect 19567 19904 19579 19907
rect 19610 19904 19616 19916
rect 19567 19876 19616 19904
rect 19567 19873 19579 19876
rect 19521 19867 19579 19873
rect 19610 19864 19616 19876
rect 19668 19864 19674 19916
rect 19429 19839 19487 19845
rect 19429 19805 19441 19839
rect 19475 19836 19487 19839
rect 19886 19836 19892 19848
rect 19475 19808 19892 19836
rect 19475 19805 19487 19808
rect 19429 19799 19487 19805
rect 19886 19796 19892 19808
rect 19944 19796 19950 19848
rect 19518 19660 19524 19712
rect 19576 19700 19582 19712
rect 19705 19703 19763 19709
rect 19705 19700 19717 19703
rect 19576 19672 19717 19700
rect 19576 19660 19582 19672
rect 19705 19669 19717 19672
rect 19751 19669 19763 19703
rect 19705 19663 19763 19669
rect 1104 19610 21712 19632
rect 1104 19558 4416 19610
rect 4468 19558 4480 19610
rect 4532 19558 4544 19610
rect 4596 19558 4608 19610
rect 4660 19558 11286 19610
rect 11338 19558 11350 19610
rect 11402 19558 11414 19610
rect 11466 19558 11478 19610
rect 11530 19558 18155 19610
rect 18207 19558 18219 19610
rect 18271 19558 18283 19610
rect 18335 19558 18347 19610
rect 18399 19558 21712 19610
rect 1104 19536 21712 19558
rect 4246 19320 4252 19372
rect 4304 19360 4310 19372
rect 5166 19360 5172 19372
rect 4304 19332 5172 19360
rect 4304 19320 4310 19332
rect 5166 19320 5172 19332
rect 5224 19320 5230 19372
rect 18874 19292 18880 19304
rect 18835 19264 18880 19292
rect 18874 19252 18880 19264
rect 18932 19252 18938 19304
rect 18966 19252 18972 19304
rect 19024 19301 19030 19304
rect 19024 19295 19047 19301
rect 19035 19261 19047 19295
rect 19024 19255 19047 19261
rect 19024 19252 19030 19255
rect 19334 19184 19340 19236
rect 19392 19224 19398 19236
rect 19429 19227 19487 19233
rect 19429 19224 19441 19227
rect 19392 19196 19441 19224
rect 19392 19184 19398 19196
rect 19429 19193 19441 19196
rect 19475 19193 19487 19227
rect 19429 19187 19487 19193
rect 1104 19066 21712 19088
rect 1104 19014 7851 19066
rect 7903 19014 7915 19066
rect 7967 19014 7979 19066
rect 8031 19014 8043 19066
rect 8095 19014 14720 19066
rect 14772 19014 14784 19066
rect 14836 19014 14848 19066
rect 14900 19014 14912 19066
rect 14964 19014 21712 19066
rect 1104 18992 21712 19014
rect 18877 18955 18935 18961
rect 18877 18921 18889 18955
rect 18923 18952 18935 18955
rect 19242 18952 19248 18964
rect 18923 18924 19248 18952
rect 18923 18921 18935 18924
rect 18877 18915 18935 18921
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 18966 18844 18972 18896
rect 19024 18884 19030 18896
rect 19024 18856 19656 18884
rect 19024 18844 19030 18856
rect 19242 18816 19248 18828
rect 19203 18788 19248 18816
rect 19242 18776 19248 18788
rect 19300 18776 19306 18828
rect 19628 18825 19656 18856
rect 19613 18819 19671 18825
rect 19613 18785 19625 18819
rect 19659 18785 19671 18819
rect 19613 18779 19671 18785
rect 19334 18748 19340 18760
rect 19295 18720 19340 18748
rect 19334 18708 19340 18720
rect 19392 18708 19398 18760
rect 19521 18751 19579 18757
rect 19521 18717 19533 18751
rect 19567 18717 19579 18751
rect 19521 18711 19579 18717
rect 18874 18640 18880 18692
rect 18932 18680 18938 18692
rect 19536 18680 19564 18711
rect 18932 18652 19564 18680
rect 18932 18640 18938 18652
rect 1104 18522 21712 18544
rect 1104 18470 4416 18522
rect 4468 18470 4480 18522
rect 4532 18470 4544 18522
rect 4596 18470 4608 18522
rect 4660 18470 11286 18522
rect 11338 18470 11350 18522
rect 11402 18470 11414 18522
rect 11466 18470 11478 18522
rect 11530 18470 18155 18522
rect 18207 18470 18219 18522
rect 18271 18470 18283 18522
rect 18335 18470 18347 18522
rect 18399 18470 21712 18522
rect 1104 18448 21712 18470
rect 18966 18272 18972 18284
rect 18800 18244 18972 18272
rect 18800 18213 18828 18244
rect 18966 18232 18972 18244
rect 19024 18232 19030 18284
rect 18785 18207 18843 18213
rect 18785 18173 18797 18207
rect 18831 18173 18843 18207
rect 18785 18167 18843 18173
rect 18800 18136 18828 18167
rect 18874 18164 18880 18216
rect 18932 18204 18938 18216
rect 19245 18207 19303 18213
rect 19245 18204 19257 18207
rect 18932 18176 19257 18204
rect 18932 18164 18938 18176
rect 19245 18173 19257 18176
rect 19291 18173 19303 18207
rect 19245 18167 19303 18173
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 19352 18136 19380 18167
rect 18800 18108 19380 18136
rect 19794 18068 19800 18080
rect 19755 18040 19800 18068
rect 19794 18028 19800 18040
rect 19852 18028 19858 18080
rect 1104 17978 21712 18000
rect 1104 17926 7851 17978
rect 7903 17926 7915 17978
rect 7967 17926 7979 17978
rect 8031 17926 8043 17978
rect 8095 17926 14720 17978
rect 14772 17926 14784 17978
rect 14836 17926 14848 17978
rect 14900 17926 14912 17978
rect 14964 17926 21712 17978
rect 1104 17904 21712 17926
rect 19886 17796 19892 17808
rect 18616 17768 19564 17796
rect 19847 17768 19892 17796
rect 18616 17737 18644 17768
rect 18601 17731 18659 17737
rect 18601 17697 18613 17731
rect 18647 17697 18659 17731
rect 18601 17691 18659 17697
rect 18785 17731 18843 17737
rect 18785 17697 18797 17731
rect 18831 17728 18843 17731
rect 19334 17728 19340 17740
rect 18831 17700 19340 17728
rect 18831 17697 18843 17700
rect 18785 17691 18843 17697
rect 19334 17688 19340 17700
rect 19392 17688 19398 17740
rect 19536 17737 19564 17768
rect 19886 17756 19892 17768
rect 19944 17756 19950 17808
rect 19521 17731 19579 17737
rect 19521 17697 19533 17731
rect 19567 17728 19579 17731
rect 19794 17728 19800 17740
rect 19567 17700 19800 17728
rect 19567 17697 19579 17700
rect 19521 17691 19579 17697
rect 19794 17688 19800 17700
rect 19852 17688 19858 17740
rect 1104 17434 21712 17456
rect 1104 17382 4416 17434
rect 4468 17382 4480 17434
rect 4532 17382 4544 17434
rect 4596 17382 4608 17434
rect 4660 17382 11286 17434
rect 11338 17382 11350 17434
rect 11402 17382 11414 17434
rect 11466 17382 11478 17434
rect 11530 17382 18155 17434
rect 18207 17382 18219 17434
rect 18271 17382 18283 17434
rect 18335 17382 18347 17434
rect 18399 17382 21712 17434
rect 1104 17360 21712 17382
rect 19334 17280 19340 17332
rect 19392 17320 19398 17332
rect 19429 17323 19487 17329
rect 19429 17320 19441 17323
rect 19392 17292 19441 17320
rect 19392 17280 19398 17292
rect 19429 17289 19441 17292
rect 19475 17289 19487 17323
rect 19429 17283 19487 17289
rect 19242 17116 19248 17128
rect 19203 17088 19248 17116
rect 19242 17076 19248 17088
rect 19300 17076 19306 17128
rect 1104 16890 21712 16912
rect 1104 16838 7851 16890
rect 7903 16838 7915 16890
rect 7967 16838 7979 16890
rect 8031 16838 8043 16890
rect 8095 16838 14720 16890
rect 14772 16838 14784 16890
rect 14836 16838 14848 16890
rect 14900 16838 14912 16890
rect 14964 16838 21712 16890
rect 1104 16816 21712 16838
rect 16393 16779 16451 16785
rect 16393 16745 16405 16779
rect 16439 16776 16451 16779
rect 17770 16776 17776 16788
rect 16439 16748 17776 16776
rect 16439 16745 16451 16748
rect 16393 16739 16451 16745
rect 17770 16736 17776 16748
rect 17828 16736 17834 16788
rect 16209 16643 16267 16649
rect 16209 16609 16221 16643
rect 16255 16640 16267 16643
rect 17862 16640 17868 16652
rect 16255 16612 17868 16640
rect 16255 16609 16267 16612
rect 16209 16603 16267 16609
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 1104 16346 21712 16368
rect 1104 16294 4416 16346
rect 4468 16294 4480 16346
rect 4532 16294 4544 16346
rect 4596 16294 4608 16346
rect 4660 16294 11286 16346
rect 11338 16294 11350 16346
rect 11402 16294 11414 16346
rect 11466 16294 11478 16346
rect 11530 16294 18155 16346
rect 18207 16294 18219 16346
rect 18271 16294 18283 16346
rect 18335 16294 18347 16346
rect 18399 16294 21712 16346
rect 1104 16272 21712 16294
rect 15749 16235 15807 16241
rect 15749 16201 15761 16235
rect 15795 16232 15807 16235
rect 19242 16232 19248 16244
rect 15795 16204 19248 16232
rect 15795 16201 15807 16204
rect 15749 16195 15807 16201
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 16206 16096 16212 16108
rect 16167 16068 16212 16096
rect 16206 16056 16212 16068
rect 16264 16056 16270 16108
rect 16390 16096 16396 16108
rect 16351 16068 16396 16096
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 16114 16028 16120 16040
rect 16075 16000 16120 16028
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 16482 16028 16488 16040
rect 16443 16000 16488 16028
rect 16482 15988 16488 16000
rect 16540 15988 16546 16040
rect 1104 15802 21712 15824
rect 1104 15750 7851 15802
rect 7903 15750 7915 15802
rect 7967 15750 7979 15802
rect 8031 15750 8043 15802
rect 8095 15750 14720 15802
rect 14772 15750 14784 15802
rect 14836 15750 14848 15802
rect 14900 15750 14912 15802
rect 14964 15750 21712 15802
rect 1104 15728 21712 15750
rect 16390 15648 16396 15700
rect 16448 15648 16454 15700
rect 17862 15648 17868 15700
rect 17920 15688 17926 15700
rect 19061 15691 19119 15697
rect 19061 15688 19073 15691
rect 17920 15660 19073 15688
rect 17920 15648 17926 15660
rect 19061 15657 19073 15660
rect 19107 15657 19119 15691
rect 19061 15651 19119 15657
rect 15838 15580 15844 15632
rect 15896 15620 15902 15632
rect 16408 15620 16436 15648
rect 15896 15592 16528 15620
rect 15896 15580 15902 15592
rect 15749 15555 15807 15561
rect 15749 15521 15761 15555
rect 15795 15552 15807 15555
rect 15930 15552 15936 15564
rect 15795 15524 15936 15552
rect 15795 15521 15807 15524
rect 15749 15515 15807 15521
rect 15930 15512 15936 15524
rect 15988 15552 15994 15564
rect 16301 15555 16359 15561
rect 16301 15552 16313 15555
rect 15988 15524 16313 15552
rect 15988 15512 15994 15524
rect 16301 15521 16313 15524
rect 16347 15552 16359 15555
rect 16390 15552 16396 15564
rect 16347 15524 16396 15552
rect 16347 15521 16359 15524
rect 16301 15515 16359 15521
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 16500 15561 16528 15592
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15521 16543 15555
rect 17770 15552 17776 15564
rect 17731 15524 17776 15552
rect 16485 15515 16543 15521
rect 17770 15512 17776 15524
rect 17828 15512 17834 15564
rect 18877 15555 18935 15561
rect 18877 15521 18889 15555
rect 18923 15521 18935 15555
rect 18877 15515 18935 15521
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15484 15715 15487
rect 15838 15484 15844 15496
rect 15703 15456 15844 15484
rect 15703 15453 15715 15456
rect 15657 15447 15715 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 18892 15484 18920 15515
rect 16684 15456 18920 15484
rect 16114 15308 16120 15360
rect 16172 15348 16178 15360
rect 16684 15348 16712 15456
rect 16172 15320 16712 15348
rect 16761 15351 16819 15357
rect 16172 15308 16178 15320
rect 16761 15317 16773 15351
rect 16807 15348 16819 15351
rect 16942 15348 16948 15360
rect 16807 15320 16948 15348
rect 16807 15317 16819 15320
rect 16761 15311 16819 15317
rect 16942 15308 16948 15320
rect 17000 15308 17006 15360
rect 17034 15308 17040 15360
rect 17092 15348 17098 15360
rect 17957 15351 18015 15357
rect 17957 15348 17969 15351
rect 17092 15320 17969 15348
rect 17092 15308 17098 15320
rect 17957 15317 17969 15320
rect 18003 15317 18015 15351
rect 17957 15311 18015 15317
rect 1104 15258 21712 15280
rect 1104 15206 4416 15258
rect 4468 15206 4480 15258
rect 4532 15206 4544 15258
rect 4596 15206 4608 15258
rect 4660 15206 11286 15258
rect 11338 15206 11350 15258
rect 11402 15206 11414 15258
rect 11466 15206 11478 15258
rect 11530 15206 18155 15258
rect 18207 15206 18219 15258
rect 18271 15206 18283 15258
rect 18335 15206 18347 15258
rect 18399 15206 21712 15258
rect 1104 15184 21712 15206
rect 16117 15147 16175 15153
rect 16117 15113 16129 15147
rect 16163 15144 16175 15147
rect 16206 15144 16212 15156
rect 16163 15116 16212 15144
rect 16163 15113 16175 15116
rect 16117 15107 16175 15113
rect 16206 15104 16212 15116
rect 16264 15104 16270 15156
rect 15838 14940 15844 14952
rect 15799 14912 15844 14940
rect 15838 14900 15844 14912
rect 15896 14900 15902 14952
rect 15930 14900 15936 14952
rect 15988 14940 15994 14952
rect 15988 14912 16033 14940
rect 15988 14900 15994 14912
rect 1104 14714 21712 14736
rect 1104 14662 7851 14714
rect 7903 14662 7915 14714
rect 7967 14662 7979 14714
rect 8031 14662 8043 14714
rect 8095 14662 14720 14714
rect 14772 14662 14784 14714
rect 14836 14662 14848 14714
rect 14900 14662 14912 14714
rect 14964 14662 21712 14714
rect 1104 14640 21712 14662
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 17034 14600 17040 14612
rect 16632 14572 17040 14600
rect 16632 14560 16638 14572
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 17589 14535 17647 14541
rect 17589 14501 17601 14535
rect 17635 14532 17647 14535
rect 18506 14532 18512 14544
rect 17635 14504 18512 14532
rect 17635 14501 17647 14504
rect 17589 14495 17647 14501
rect 18506 14492 18512 14504
rect 18564 14492 18570 14544
rect 13357 14467 13415 14473
rect 13357 14433 13369 14467
rect 13403 14464 13415 14467
rect 14550 14464 14556 14476
rect 13403 14436 14556 14464
rect 13403 14433 13415 14436
rect 13357 14427 13415 14433
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 16485 14467 16543 14473
rect 16485 14433 16497 14467
rect 16531 14464 16543 14467
rect 16574 14464 16580 14476
rect 16531 14436 16580 14464
rect 16531 14433 16543 14436
rect 16485 14427 16543 14433
rect 16574 14424 16580 14436
rect 16632 14424 16638 14476
rect 16942 14464 16948 14476
rect 16684 14436 16948 14464
rect 16393 14399 16451 14405
rect 16393 14365 16405 14399
rect 16439 14396 16451 14399
rect 16684 14396 16712 14436
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 17034 14424 17040 14476
rect 17092 14464 17098 14476
rect 17092 14436 17137 14464
rect 17092 14424 17098 14436
rect 16439 14368 16712 14396
rect 16439 14365 16451 14368
rect 16393 14359 16451 14365
rect 13541 14263 13599 14269
rect 13541 14229 13553 14263
rect 13587 14260 13599 14263
rect 14366 14260 14372 14272
rect 13587 14232 14372 14260
rect 13587 14229 13599 14232
rect 13541 14223 13599 14229
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 1104 14170 21712 14192
rect 1104 14118 4416 14170
rect 4468 14118 4480 14170
rect 4532 14118 4544 14170
rect 4596 14118 4608 14170
rect 4660 14118 11286 14170
rect 11338 14118 11350 14170
rect 11402 14118 11414 14170
rect 11466 14118 11478 14170
rect 11530 14118 18155 14170
rect 18207 14118 18219 14170
rect 18271 14118 18283 14170
rect 18335 14118 18347 14170
rect 18399 14118 21712 14170
rect 1104 14096 21712 14118
rect 14550 14056 14556 14068
rect 14511 14028 14556 14056
rect 14550 14016 14556 14028
rect 14608 14016 14614 14068
rect 12434 13880 12440 13932
rect 12492 13920 12498 13932
rect 12492 13892 13124 13920
rect 12492 13880 12498 13892
rect 13096 13861 13124 13892
rect 12989 13855 13047 13861
rect 12989 13821 13001 13855
rect 13035 13821 13047 13855
rect 12989 13815 13047 13821
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13852 13139 13855
rect 13446 13852 13452 13864
rect 13127 13824 13452 13852
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 13004 13716 13032 13815
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 14369 13855 14427 13861
rect 14369 13852 14381 13855
rect 13688 13824 14381 13852
rect 13688 13812 13694 13824
rect 14369 13821 14381 13824
rect 14415 13821 14427 13855
rect 14369 13815 14427 13821
rect 13354 13744 13360 13796
rect 13412 13784 13418 13796
rect 13541 13787 13599 13793
rect 13541 13784 13553 13787
rect 13412 13756 13553 13784
rect 13412 13744 13418 13756
rect 13541 13753 13553 13756
rect 13587 13753 13599 13787
rect 13541 13747 13599 13753
rect 13722 13716 13728 13728
rect 13004 13688 13728 13716
rect 13722 13676 13728 13688
rect 13780 13676 13786 13728
rect 1104 13626 21712 13648
rect 1104 13574 7851 13626
rect 7903 13574 7915 13626
rect 7967 13574 7979 13626
rect 8031 13574 8043 13626
rect 8095 13574 14720 13626
rect 14772 13574 14784 13626
rect 14836 13574 14848 13626
rect 14900 13574 14912 13626
rect 14964 13574 21712 13626
rect 1104 13552 21712 13574
rect 12897 13515 12955 13521
rect 12897 13481 12909 13515
rect 12943 13512 12955 13515
rect 16114 13512 16120 13524
rect 12943 13484 16120 13512
rect 12943 13481 12955 13484
rect 12897 13475 12955 13481
rect 16114 13472 16120 13484
rect 16172 13472 16178 13524
rect 13262 13376 13268 13388
rect 13223 13348 13268 13376
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 13446 13336 13452 13388
rect 13504 13376 13510 13388
rect 13633 13379 13691 13385
rect 13633 13376 13645 13379
rect 13504 13348 13645 13376
rect 13504 13336 13510 13348
rect 13633 13345 13645 13348
rect 13679 13345 13691 13379
rect 13633 13339 13691 13345
rect 13722 13336 13728 13388
rect 13780 13376 13786 13388
rect 13780 13348 13825 13376
rect 13780 13336 13786 13348
rect 13354 13308 13360 13320
rect 13315 13280 13360 13308
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 1104 13082 21712 13104
rect 1104 13030 4416 13082
rect 4468 13030 4480 13082
rect 4532 13030 4544 13082
rect 4596 13030 4608 13082
rect 4660 13030 11286 13082
rect 11338 13030 11350 13082
rect 11402 13030 11414 13082
rect 11466 13030 11478 13082
rect 11530 13030 18155 13082
rect 18207 13030 18219 13082
rect 18271 13030 18283 13082
rect 18335 13030 18347 13082
rect 18399 13030 21712 13082
rect 1104 13008 21712 13030
rect 13538 12724 13544 12776
rect 13596 12764 13602 12776
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 13596 12736 13645 12764
rect 13596 12724 13602 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 13725 12767 13783 12773
rect 13725 12733 13737 12767
rect 13771 12764 13783 12767
rect 13998 12764 14004 12776
rect 13771 12736 14004 12764
rect 13771 12733 13783 12736
rect 13725 12727 13783 12733
rect 13648 12696 13676 12727
rect 13998 12724 14004 12736
rect 14056 12764 14062 12776
rect 14093 12767 14151 12773
rect 14093 12764 14105 12767
rect 14056 12736 14105 12764
rect 14056 12724 14062 12736
rect 14093 12733 14105 12736
rect 14139 12733 14151 12767
rect 14093 12727 14151 12733
rect 14185 12767 14243 12773
rect 14185 12733 14197 12767
rect 14231 12733 14243 12767
rect 14185 12727 14243 12733
rect 14200 12696 14228 12727
rect 14366 12724 14372 12776
rect 14424 12764 14430 12776
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 14424 12736 15669 12764
rect 14424 12724 14430 12736
rect 15657 12733 15669 12736
rect 15703 12733 15715 12767
rect 15657 12727 15715 12733
rect 13648 12668 14228 12696
rect 14737 12699 14795 12705
rect 14737 12665 14749 12699
rect 14783 12696 14795 12699
rect 19150 12696 19156 12708
rect 14783 12668 19156 12696
rect 14783 12665 14795 12668
rect 14737 12659 14795 12665
rect 19150 12656 19156 12668
rect 19208 12656 19214 12708
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 15841 12631 15899 12637
rect 15841 12628 15853 12631
rect 13872 12600 15853 12628
rect 13872 12588 13878 12600
rect 15841 12597 15853 12600
rect 15887 12597 15899 12631
rect 15841 12591 15899 12597
rect 1104 12538 21712 12560
rect 1104 12486 7851 12538
rect 7903 12486 7915 12538
rect 7967 12486 7979 12538
rect 8031 12486 8043 12538
rect 8095 12486 14720 12538
rect 14772 12486 14784 12538
rect 14836 12486 14848 12538
rect 14900 12486 14912 12538
rect 14964 12486 21712 12538
rect 1104 12464 21712 12486
rect 13722 12356 13728 12368
rect 12728 12328 13728 12356
rect 12728 12232 12756 12328
rect 12897 12291 12955 12297
rect 12897 12257 12909 12291
rect 12943 12288 12955 12291
rect 13446 12288 13452 12300
rect 12943 12260 13452 12288
rect 12943 12257 12955 12260
rect 12897 12251 12955 12257
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 13648 12297 13676 12328
rect 13722 12316 13728 12328
rect 13780 12316 13786 12368
rect 13998 12356 14004 12368
rect 13959 12328 14004 12356
rect 13998 12316 14004 12328
rect 14056 12316 14062 12368
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12257 13691 12291
rect 13633 12251 13691 12257
rect 12710 12220 12716 12232
rect 12671 12192 12716 12220
rect 12710 12180 12716 12192
rect 12768 12180 12774 12232
rect 1104 11994 21712 12016
rect 1104 11942 4416 11994
rect 4468 11942 4480 11994
rect 4532 11942 4544 11994
rect 4596 11942 4608 11994
rect 4660 11942 11286 11994
rect 11338 11942 11350 11994
rect 11402 11942 11414 11994
rect 11466 11942 11478 11994
rect 11530 11942 18155 11994
rect 18207 11942 18219 11994
rect 18271 11942 18283 11994
rect 18335 11942 18347 11994
rect 18399 11942 21712 11994
rect 1104 11920 21712 11942
rect 13538 11880 13544 11892
rect 13499 11852 13544 11880
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 10502 11676 10508 11688
rect 10463 11648 10508 11676
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 13357 11679 13415 11685
rect 13357 11645 13369 11679
rect 13403 11676 13415 11679
rect 13814 11676 13820 11688
rect 13403 11648 13820 11676
rect 13403 11645 13415 11648
rect 13357 11639 13415 11645
rect 13814 11636 13820 11648
rect 13872 11636 13878 11688
rect 10689 11543 10747 11549
rect 10689 11509 10701 11543
rect 10735 11540 10747 11543
rect 11698 11540 11704 11552
rect 10735 11512 11704 11540
rect 10735 11509 10747 11512
rect 10689 11503 10747 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 1104 11450 21712 11472
rect 1104 11398 7851 11450
rect 7903 11398 7915 11450
rect 7967 11398 7979 11450
rect 8031 11398 8043 11450
rect 8095 11398 14720 11450
rect 14772 11398 14784 11450
rect 14836 11398 14848 11450
rect 14900 11398 14912 11450
rect 14964 11398 21712 11450
rect 1104 11376 21712 11398
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 10689 11339 10747 11345
rect 10689 11336 10701 11339
rect 10652 11308 10701 11336
rect 10652 11296 10658 11308
rect 10689 11305 10701 11308
rect 10735 11305 10747 11339
rect 10689 11299 10747 11305
rect 13541 11339 13599 11345
rect 13541 11305 13553 11339
rect 13587 11336 13599 11339
rect 13630 11336 13636 11348
rect 13587 11308 13636 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11200 10563 11203
rect 11146 11200 11152 11212
rect 10551 11172 11152 11200
rect 10551 11169 10563 11172
rect 10505 11163 10563 11169
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 11609 11203 11667 11209
rect 11609 11169 11621 11203
rect 11655 11169 11667 11203
rect 13354 11200 13360 11212
rect 13315 11172 13360 11200
rect 11609 11163 11667 11169
rect 10410 11092 10416 11144
rect 10468 11132 10474 11144
rect 11624 11132 11652 11163
rect 13354 11160 13360 11172
rect 13412 11160 13418 11212
rect 10468 11104 11652 11132
rect 10468 11092 10474 11104
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 11793 11067 11851 11073
rect 11793 11064 11805 11067
rect 9732 11036 11805 11064
rect 9732 11024 9738 11036
rect 11793 11033 11805 11036
rect 11839 11033 11851 11067
rect 11793 11027 11851 11033
rect 1104 10906 21712 10928
rect 1104 10854 4416 10906
rect 4468 10854 4480 10906
rect 4532 10854 4544 10906
rect 4596 10854 4608 10906
rect 4660 10854 11286 10906
rect 11338 10854 11350 10906
rect 11402 10854 11414 10906
rect 11466 10854 11478 10906
rect 11530 10854 18155 10906
rect 18207 10854 18219 10906
rect 18271 10854 18283 10906
rect 18335 10854 18347 10906
rect 18399 10854 21712 10906
rect 1104 10832 21712 10854
rect 9217 10795 9275 10801
rect 9217 10761 9229 10795
rect 9263 10792 9275 10795
rect 10502 10792 10508 10804
rect 9263 10764 10508 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10588 9091 10591
rect 9674 10588 9680 10600
rect 9079 10560 9680 10588
rect 9079 10557 9091 10560
rect 9033 10551 9091 10557
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 9950 10548 9956 10600
rect 10008 10588 10014 10600
rect 10137 10591 10195 10597
rect 10137 10588 10149 10591
rect 10008 10560 10149 10588
rect 10008 10548 10014 10560
rect 10137 10557 10149 10560
rect 10183 10557 10195 10591
rect 10137 10551 10195 10557
rect 10226 10548 10232 10600
rect 10284 10588 10290 10600
rect 10284 10560 10329 10588
rect 10284 10548 10290 10560
rect 10502 10480 10508 10532
rect 10560 10520 10566 10532
rect 10689 10523 10747 10529
rect 10689 10520 10701 10523
rect 10560 10492 10701 10520
rect 10560 10480 10566 10492
rect 10689 10489 10701 10492
rect 10735 10489 10747 10523
rect 10689 10483 10747 10489
rect 1104 10362 21712 10384
rect 1104 10310 7851 10362
rect 7903 10310 7915 10362
rect 7967 10310 7979 10362
rect 8031 10310 8043 10362
rect 8095 10310 14720 10362
rect 14772 10310 14784 10362
rect 14836 10310 14848 10362
rect 14900 10310 14912 10362
rect 14964 10310 21712 10362
rect 1104 10288 21712 10310
rect 11146 10208 11152 10260
rect 11204 10248 11210 10260
rect 12989 10251 13047 10257
rect 12989 10248 13001 10251
rect 11204 10220 13001 10248
rect 11204 10208 11210 10220
rect 12989 10217 13001 10220
rect 13035 10217 13047 10251
rect 12989 10211 13047 10217
rect 10796 10152 11376 10180
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 10796 10121 10824 10152
rect 10781 10115 10839 10121
rect 10781 10112 10793 10115
rect 10744 10084 10793 10112
rect 10744 10072 10750 10084
rect 10781 10081 10793 10084
rect 10827 10081 10839 10115
rect 10781 10075 10839 10081
rect 10873 10115 10931 10121
rect 10873 10081 10885 10115
rect 10919 10112 10931 10115
rect 11146 10112 11152 10124
rect 10919 10084 11152 10112
rect 10919 10081 10931 10084
rect 10873 10075 10931 10081
rect 11146 10072 11152 10084
rect 11204 10112 11210 10124
rect 11348 10121 11376 10152
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 11204 10084 11253 10112
rect 11204 10072 11210 10084
rect 11241 10081 11253 10084
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 11333 10115 11391 10121
rect 11333 10081 11345 10115
rect 11379 10081 11391 10115
rect 11333 10075 11391 10081
rect 11698 10072 11704 10124
rect 11756 10112 11762 10124
rect 12805 10115 12863 10121
rect 12805 10112 12817 10115
rect 11756 10084 12817 10112
rect 11756 10072 11762 10084
rect 12805 10081 12817 10084
rect 12851 10081 12863 10115
rect 12805 10075 12863 10081
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 19242 10044 19248 10056
rect 11931 10016 19248 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 1104 9818 21712 9840
rect 1104 9766 4416 9818
rect 4468 9766 4480 9818
rect 4532 9766 4544 9818
rect 4596 9766 4608 9818
rect 4660 9766 11286 9818
rect 11338 9766 11350 9818
rect 11402 9766 11414 9818
rect 11466 9766 11478 9818
rect 11530 9766 18155 9818
rect 18207 9766 18219 9818
rect 18271 9766 18283 9818
rect 18335 9766 18347 9818
rect 18399 9766 21712 9818
rect 1104 9744 21712 9766
rect 11057 9707 11115 9713
rect 11057 9673 11069 9707
rect 11103 9704 11115 9707
rect 11146 9704 11152 9716
rect 11103 9676 11152 9704
rect 11103 9673 11115 9676
rect 11057 9667 11115 9673
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 5166 9596 5172 9648
rect 5224 9636 5230 9648
rect 5350 9636 5356 9648
rect 5224 9608 5356 9636
rect 5224 9596 5230 9608
rect 5350 9596 5356 9608
rect 5408 9596 5414 9648
rect 9950 9568 9956 9580
rect 9911 9540 9956 9568
rect 9950 9528 9956 9540
rect 10008 9568 10014 9580
rect 10008 9540 10272 9568
rect 10008 9528 10014 9540
rect 10045 9503 10103 9509
rect 10045 9469 10057 9503
rect 10091 9500 10103 9503
rect 10134 9500 10140 9512
rect 10091 9472 10140 9500
rect 10091 9469 10103 9472
rect 10045 9463 10103 9469
rect 10134 9460 10140 9472
rect 10192 9460 10198 9512
rect 10244 9500 10272 9540
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 10244 9472 10517 9500
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 10505 9463 10563 9469
rect 10597 9503 10655 9509
rect 10597 9469 10609 9503
rect 10643 9469 10655 9503
rect 10597 9463 10655 9469
rect 10152 9432 10180 9460
rect 10612 9432 10640 9463
rect 10778 9432 10784 9444
rect 10152 9404 10784 9432
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 1104 9274 21712 9296
rect 1104 9222 7851 9274
rect 7903 9222 7915 9274
rect 7967 9222 7979 9274
rect 8031 9222 8043 9274
rect 8095 9222 14720 9274
rect 14772 9222 14784 9274
rect 14836 9222 14848 9274
rect 14900 9222 14912 9274
rect 14964 9222 21712 9274
rect 1104 9200 21712 9222
rect 10045 9163 10103 9169
rect 10045 9129 10057 9163
rect 10091 9160 10103 9163
rect 13354 9160 13360 9172
rect 10091 9132 13360 9160
rect 10091 9129 10103 9132
rect 10045 9123 10103 9129
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 7650 9024 7656 9036
rect 7611 8996 7656 9024
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 10410 9024 10416 9036
rect 10371 8996 10416 9024
rect 10410 8984 10416 8996
rect 10468 8984 10474 9036
rect 10778 9024 10784 9036
rect 10739 8996 10784 9024
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 10502 8956 10508 8968
rect 10463 8928 10508 8956
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8925 10747 8959
rect 10689 8919 10747 8925
rect 9950 8848 9956 8900
rect 10008 8888 10014 8900
rect 10704 8888 10732 8919
rect 10008 8860 10732 8888
rect 10008 8848 10014 8860
rect 7837 8823 7895 8829
rect 7837 8789 7849 8823
rect 7883 8820 7895 8823
rect 9582 8820 9588 8832
rect 7883 8792 9588 8820
rect 7883 8789 7895 8792
rect 7837 8783 7895 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 1104 8730 21712 8752
rect 1104 8678 4416 8730
rect 4468 8678 4480 8730
rect 4532 8678 4544 8730
rect 4596 8678 4608 8730
rect 4660 8678 11286 8730
rect 11338 8678 11350 8730
rect 11402 8678 11414 8730
rect 11466 8678 11478 8730
rect 11530 8678 18155 8730
rect 18207 8678 18219 8730
rect 18271 8678 18283 8730
rect 18335 8678 18347 8730
rect 18399 8678 21712 8730
rect 1104 8656 21712 8678
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 7837 8619 7895 8625
rect 7837 8616 7849 8619
rect 5960 8588 7849 8616
rect 5960 8576 5966 8588
rect 7837 8585 7849 8588
rect 7883 8585 7895 8619
rect 10686 8616 10692 8628
rect 10647 8588 10692 8616
rect 7837 8579 7895 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 2409 8551 2467 8557
rect 2409 8517 2421 8551
rect 2455 8548 2467 8551
rect 3050 8548 3056 8560
rect 2455 8520 3056 8548
rect 2455 8517 2467 8520
rect 2409 8511 2467 8517
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 6914 8508 6920 8560
rect 6972 8548 6978 8560
rect 8941 8551 8999 8557
rect 8941 8548 8953 8551
rect 6972 8520 8953 8548
rect 6972 8508 6978 8520
rect 8941 8517 8953 8520
rect 8987 8517 8999 8551
rect 8941 8511 8999 8517
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8412 2283 8415
rect 2590 8412 2596 8424
rect 2271 8384 2596 8412
rect 2271 8381 2283 8384
rect 2225 8375 2283 8381
rect 2590 8372 2596 8384
rect 2648 8372 2654 8424
rect 7653 8415 7711 8421
rect 7653 8381 7665 8415
rect 7699 8412 7711 8415
rect 8662 8412 8668 8424
rect 7699 8384 8668 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 10505 8415 10563 8421
rect 8812 8384 8857 8412
rect 8812 8372 8818 8384
rect 10505 8381 10517 8415
rect 10551 8412 10563 8415
rect 10594 8412 10600 8424
rect 10551 8384 10600 8412
rect 10551 8381 10563 8384
rect 10505 8375 10563 8381
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 1104 8186 21712 8208
rect 1104 8134 7851 8186
rect 7903 8134 7915 8186
rect 7967 8134 7979 8186
rect 8031 8134 8043 8186
rect 8095 8134 14720 8186
rect 14772 8134 14784 8186
rect 14836 8134 14848 8186
rect 14900 8134 14912 8186
rect 14964 8134 21712 8186
rect 1104 8112 21712 8134
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 7650 8072 7656 8084
rect 6411 8044 7656 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7936 2283 7939
rect 2498 7936 2504 7948
rect 2271 7908 2504 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 4706 7896 4712 7948
rect 4764 7936 4770 7948
rect 4801 7939 4859 7945
rect 4801 7936 4813 7939
rect 4764 7908 4813 7936
rect 4764 7896 4770 7908
rect 4801 7905 4813 7908
rect 4847 7905 4859 7939
rect 4801 7899 4859 7905
rect 6181 7939 6239 7945
rect 6181 7905 6193 7939
rect 6227 7936 6239 7939
rect 6914 7936 6920 7948
rect 6227 7908 6920 7936
rect 6227 7905 6239 7908
rect 6181 7899 6239 7905
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 7156 7908 7389 7936
rect 7156 7896 7162 7908
rect 7377 7905 7389 7908
rect 7423 7905 7435 7939
rect 7377 7899 7435 7905
rect 7282 7868 7288 7880
rect 7243 7840 7288 7868
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 2314 7692 2320 7744
rect 2372 7732 2378 7744
rect 2409 7735 2467 7741
rect 2409 7732 2421 7735
rect 2372 7704 2421 7732
rect 2372 7692 2378 7704
rect 2409 7701 2421 7704
rect 2455 7701 2467 7735
rect 2409 7695 2467 7701
rect 4985 7735 5043 7741
rect 4985 7701 4997 7735
rect 5031 7732 5043 7735
rect 6822 7732 6828 7744
rect 5031 7704 6828 7732
rect 5031 7701 5043 7704
rect 4985 7695 5043 7701
rect 6822 7692 6828 7704
rect 6880 7692 6886 7744
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 7524 7704 7573 7732
rect 7524 7692 7530 7704
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 1104 7642 21712 7664
rect 1104 7590 4416 7642
rect 4468 7590 4480 7642
rect 4532 7590 4544 7642
rect 4596 7590 4608 7642
rect 4660 7590 11286 7642
rect 11338 7590 11350 7642
rect 11402 7590 11414 7642
rect 11466 7590 11478 7642
rect 11530 7590 18155 7642
rect 18207 7590 18219 7642
rect 18271 7590 18283 7642
rect 18335 7590 18347 7642
rect 18399 7590 21712 7642
rect 1104 7568 21712 7590
rect 8662 7488 8668 7540
rect 8720 7528 8726 7540
rect 10045 7531 10103 7537
rect 10045 7528 10057 7531
rect 8720 7500 10057 7528
rect 8720 7488 8726 7500
rect 10045 7497 10057 7500
rect 10091 7497 10103 7531
rect 10045 7491 10103 7497
rect 7742 7392 7748 7404
rect 7703 7364 7748 7392
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 2406 7324 2412 7336
rect 2271 7296 2412 7324
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 3329 7327 3387 7333
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 3510 7324 3516 7336
rect 3375 7296 3516 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 3510 7284 3516 7296
rect 3568 7284 3574 7336
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7324 4859 7327
rect 4982 7324 4988 7336
rect 4847 7296 4988 7324
rect 4847 7293 4859 7296
rect 4801 7287 4859 7293
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 7837 7327 7895 7333
rect 7837 7293 7849 7327
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 7852 7256 7880 7287
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 8297 7327 8355 7333
rect 8297 7324 8309 7327
rect 8260 7296 8309 7324
rect 8260 7284 8266 7296
rect 8297 7293 8309 7296
rect 8343 7293 8355 7327
rect 8297 7287 8355 7293
rect 8389 7327 8447 7333
rect 8389 7293 8401 7327
rect 8435 7293 8447 7327
rect 8389 7287 8447 7293
rect 8220 7256 8248 7284
rect 7852 7228 8248 7256
rect 2222 7148 2228 7200
rect 2280 7188 2286 7200
rect 2409 7191 2467 7197
rect 2409 7188 2421 7191
rect 2280 7160 2421 7188
rect 2280 7148 2286 7160
rect 2409 7157 2421 7160
rect 2455 7157 2467 7191
rect 2409 7151 2467 7157
rect 3142 7148 3148 7200
rect 3200 7188 3206 7200
rect 3513 7191 3571 7197
rect 3513 7188 3525 7191
rect 3200 7160 3525 7188
rect 3200 7148 3206 7160
rect 3513 7157 3525 7160
rect 3559 7157 3571 7191
rect 3513 7151 3571 7157
rect 4798 7148 4804 7200
rect 4856 7188 4862 7200
rect 4985 7191 5043 7197
rect 4985 7188 4997 7191
rect 4856 7160 4997 7188
rect 4856 7148 4862 7160
rect 4985 7157 4997 7160
rect 5031 7157 5043 7191
rect 4985 7151 5043 7157
rect 7742 7148 7748 7200
rect 7800 7188 7806 7200
rect 8404 7188 8432 7287
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 9861 7327 9919 7333
rect 9861 7324 9873 7327
rect 9640 7296 9873 7324
rect 9640 7284 9646 7296
rect 9861 7293 9873 7296
rect 9907 7293 9919 7327
rect 9861 7287 9919 7293
rect 8846 7188 8852 7200
rect 7800 7160 8432 7188
rect 8807 7160 8852 7188
rect 7800 7148 7806 7160
rect 8846 7148 8852 7160
rect 8904 7148 8910 7200
rect 1104 7098 21712 7120
rect 1104 7046 7851 7098
rect 7903 7046 7915 7098
rect 7967 7046 7979 7098
rect 8031 7046 8043 7098
rect 8095 7046 14720 7098
rect 14772 7046 14784 7098
rect 14836 7046 14848 7098
rect 14900 7046 14912 7098
rect 14964 7046 21712 7098
rect 1104 7024 21712 7046
rect 8202 6984 8208 6996
rect 8163 6956 8208 6984
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 8846 6944 8852 6996
rect 8904 6984 8910 6996
rect 18046 6984 18052 6996
rect 8904 6956 18052 6984
rect 8904 6944 8910 6956
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 7282 6876 7288 6928
rect 7340 6916 7346 6928
rect 7834 6916 7840 6928
rect 7340 6888 7840 6916
rect 7340 6876 7346 6888
rect 7834 6876 7840 6888
rect 7892 6916 7898 6928
rect 7892 6888 7972 6916
rect 7892 6876 7898 6888
rect 2222 6848 2228 6860
rect 2183 6820 2228 6848
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 4798 6848 4804 6860
rect 4759 6820 4804 6848
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 5902 6848 5908 6860
rect 5863 6820 5908 6848
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 7944 6857 7972 6888
rect 7193 6851 7251 6857
rect 7193 6848 7205 6851
rect 7156 6820 7205 6848
rect 7156 6808 7162 6820
rect 7193 6817 7205 6820
rect 7239 6848 7251 6851
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 7239 6820 7757 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 7745 6811 7803 6817
rect 7929 6851 7987 6857
rect 7929 6817 7941 6851
rect 7975 6817 7987 6851
rect 7929 6811 7987 6817
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 7282 6780 7288 6792
rect 7055 6752 7288 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 3326 6644 3332 6656
rect 2455 6616 3332 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 4890 6604 4896 6656
rect 4948 6644 4954 6656
rect 4985 6647 5043 6653
rect 4985 6644 4997 6647
rect 4948 6616 4997 6644
rect 4948 6604 4954 6616
rect 4985 6613 4997 6616
rect 5031 6613 5043 6647
rect 4985 6607 5043 6613
rect 6089 6647 6147 6653
rect 6089 6613 6101 6647
rect 6135 6644 6147 6647
rect 7650 6644 7656 6656
rect 6135 6616 7656 6644
rect 6135 6613 6147 6616
rect 6089 6607 6147 6613
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 1104 6554 21712 6576
rect 1104 6502 4416 6554
rect 4468 6502 4480 6554
rect 4532 6502 4544 6554
rect 4596 6502 4608 6554
rect 4660 6502 11286 6554
rect 11338 6502 11350 6554
rect 11402 6502 11414 6554
rect 11466 6502 11478 6554
rect 11530 6502 18155 6554
rect 18207 6502 18219 6554
rect 18271 6502 18283 6554
rect 18335 6502 18347 6554
rect 18399 6502 21712 6554
rect 1104 6480 21712 6502
rect 7193 6443 7251 6449
rect 7193 6409 7205 6443
rect 7239 6440 7251 6443
rect 10410 6440 10416 6452
rect 7239 6412 10416 6440
rect 7239 6409 7251 6412
rect 7193 6403 7251 6409
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 4246 6332 4252 6384
rect 4304 6372 4310 6384
rect 8754 6372 8760 6384
rect 4304 6344 4936 6372
rect 4304 6332 4310 6344
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6304 1823 6307
rect 2130 6304 2136 6316
rect 1811 6276 2136 6304
rect 1811 6273 1823 6276
rect 1765 6267 1823 6273
rect 2130 6264 2136 6276
rect 2188 6304 2194 6316
rect 2682 6304 2688 6316
rect 2188 6276 2688 6304
rect 2188 6264 2194 6276
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 4798 6304 4804 6316
rect 4759 6276 4804 6304
rect 4798 6264 4804 6276
rect 4856 6264 4862 6316
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 1946 6236 1952 6248
rect 1903 6208 1952 6236
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 1946 6196 1952 6208
rect 2004 6196 2010 6248
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6205 4767 6239
rect 4908 6236 4936 6344
rect 7576 6344 8760 6372
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 5031 6239 5089 6245
rect 5031 6236 5043 6239
rect 4908 6208 5043 6236
rect 4709 6199 4767 6205
rect 5031 6205 5043 6208
rect 5077 6205 5089 6239
rect 5031 6199 5089 6205
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6236 5319 6239
rect 5350 6236 5356 6248
rect 5307 6208 5356 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 2222 6128 2228 6180
rect 2280 6168 2286 6180
rect 2317 6171 2375 6177
rect 2317 6168 2329 6171
rect 2280 6140 2329 6168
rect 2280 6128 2286 6140
rect 2317 6137 2329 6140
rect 2363 6137 2375 6171
rect 4724 6168 4752 6199
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 7576 6245 7604 6344
rect 8754 6332 8760 6344
rect 8812 6332 8818 6384
rect 7834 6304 7840 6316
rect 7795 6276 7840 6304
rect 7834 6264 7840 6276
rect 7892 6264 7898 6316
rect 7561 6239 7619 6245
rect 7561 6236 7573 6239
rect 6840 6208 7573 6236
rect 5902 6168 5908 6180
rect 4724 6140 5908 6168
rect 2317 6131 2375 6137
rect 5902 6128 5908 6140
rect 5960 6128 5966 6180
rect 4341 6103 4399 6109
rect 4341 6069 4353 6103
rect 4387 6100 4399 6103
rect 6840 6100 6868 6208
rect 7561 6205 7573 6208
rect 7607 6205 7619 6239
rect 7561 6199 7619 6205
rect 7929 6239 7987 6245
rect 7929 6205 7941 6239
rect 7975 6205 7987 6239
rect 7929 6199 7987 6205
rect 7098 6128 7104 6180
rect 7156 6168 7162 6180
rect 7944 6168 7972 6199
rect 7156 6140 7972 6168
rect 7156 6128 7162 6140
rect 4387 6072 6868 6100
rect 4387 6069 4399 6072
rect 4341 6063 4399 6069
rect 1104 6010 21712 6032
rect 1104 5958 7851 6010
rect 7903 5958 7915 6010
rect 7967 5958 7979 6010
rect 8031 5958 8043 6010
rect 8095 5958 14720 6010
rect 14772 5958 14784 6010
rect 14836 5958 14848 6010
rect 14900 5958 14912 6010
rect 14964 5958 21712 6010
rect 1104 5936 21712 5958
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 7800 5868 7849 5896
rect 7800 5856 7806 5868
rect 7837 5865 7849 5868
rect 7883 5865 7895 5899
rect 7837 5859 7895 5865
rect 4908 5800 5580 5828
rect 4908 5772 4936 5800
rect 2041 5763 2099 5769
rect 2041 5729 2053 5763
rect 2087 5760 2099 5763
rect 2222 5760 2228 5772
rect 2087 5732 2228 5760
rect 2087 5729 2099 5732
rect 2041 5723 2099 5729
rect 2222 5720 2228 5732
rect 2280 5720 2286 5772
rect 2409 5763 2467 5769
rect 2409 5729 2421 5763
rect 2455 5729 2467 5763
rect 2409 5723 2467 5729
rect 2593 5763 2651 5769
rect 2593 5729 2605 5763
rect 2639 5760 2651 5763
rect 2682 5760 2688 5772
rect 2639 5732 2688 5760
rect 2639 5729 2651 5732
rect 2593 5723 2651 5729
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 1872 5624 1900 5655
rect 1946 5652 1952 5704
rect 2004 5692 2010 5704
rect 2424 5692 2452 5723
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 4801 5763 4859 5769
rect 4801 5729 4813 5763
rect 4847 5760 4859 5763
rect 4890 5760 4896 5772
rect 4847 5732 4896 5760
rect 4847 5729 4859 5732
rect 4801 5723 4859 5729
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 4985 5763 5043 5769
rect 4985 5729 4997 5763
rect 5031 5760 5043 5763
rect 5350 5760 5356 5772
rect 5031 5732 5356 5760
rect 5031 5729 5043 5732
rect 4985 5723 5043 5729
rect 5350 5720 5356 5732
rect 5408 5760 5414 5772
rect 5552 5769 5580 5800
rect 5445 5763 5503 5769
rect 5445 5760 5457 5763
rect 5408 5732 5457 5760
rect 5408 5720 5414 5732
rect 5445 5729 5457 5732
rect 5491 5729 5503 5763
rect 5445 5723 5503 5729
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5729 5595 5763
rect 7650 5760 7656 5772
rect 7611 5732 7656 5760
rect 5537 5723 5595 5729
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 2004 5664 2452 5692
rect 2004 5652 2010 5664
rect 2866 5624 2872 5636
rect 1872 5596 2872 5624
rect 2866 5584 2872 5596
rect 2924 5584 2930 5636
rect 5997 5627 6055 5633
rect 5997 5593 6009 5627
rect 6043 5624 6055 5627
rect 18782 5624 18788 5636
rect 6043 5596 18788 5624
rect 6043 5593 6055 5596
rect 5997 5587 6055 5593
rect 18782 5584 18788 5596
rect 18840 5584 18846 5636
rect 1673 5559 1731 5565
rect 1673 5525 1685 5559
rect 1719 5556 1731 5559
rect 5902 5556 5908 5568
rect 1719 5528 5908 5556
rect 1719 5525 1731 5528
rect 1673 5519 1731 5525
rect 5902 5516 5908 5528
rect 5960 5516 5966 5568
rect 1104 5466 21712 5488
rect 1104 5414 4416 5466
rect 4468 5414 4480 5466
rect 4532 5414 4544 5466
rect 4596 5414 4608 5466
rect 4660 5414 11286 5466
rect 11338 5414 11350 5466
rect 11402 5414 11414 5466
rect 11466 5414 11478 5466
rect 11530 5414 18155 5466
rect 18207 5414 18219 5466
rect 18271 5414 18283 5466
rect 18335 5414 18347 5466
rect 18399 5414 21712 5466
rect 1104 5392 21712 5414
rect 5350 5352 5356 5364
rect 5311 5324 5356 5352
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 5258 5284 5264 5296
rect 4540 5256 5264 5284
rect 2038 5216 2044 5228
rect 1999 5188 2044 5216
rect 2038 5176 2044 5188
rect 2096 5216 2102 5228
rect 2096 5188 2268 5216
rect 2096 5176 2102 5188
rect 2130 5148 2136 5160
rect 2091 5120 2136 5148
rect 2130 5108 2136 5120
rect 2188 5108 2194 5160
rect 2240 5148 2268 5188
rect 2593 5151 2651 5157
rect 2593 5148 2605 5151
rect 2240 5120 2605 5148
rect 2593 5117 2605 5120
rect 2639 5117 2651 5151
rect 2593 5111 2651 5117
rect 2685 5151 2743 5157
rect 2685 5117 2697 5151
rect 2731 5117 2743 5151
rect 2685 5111 2743 5117
rect 2148 5080 2176 5108
rect 2700 5080 2728 5111
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 4304 5120 4353 5148
rect 4304 5108 4310 5120
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 2148 5052 2728 5080
rect 3237 5083 3295 5089
rect 3237 5049 3249 5083
rect 3283 5080 3295 5083
rect 4062 5080 4068 5092
rect 3283 5052 4068 5080
rect 3283 5049 3295 5052
rect 3237 5043 3295 5049
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 4356 5080 4384 5111
rect 4430 5108 4436 5160
rect 4488 5148 4494 5160
rect 4540 5148 4568 5256
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 4893 5151 4951 5157
rect 4488 5120 4581 5148
rect 4488 5108 4494 5120
rect 4893 5117 4905 5151
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5148 5135 5151
rect 5258 5148 5264 5160
rect 5123 5120 5264 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 4908 5080 4936 5111
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 6822 5148 6828 5160
rect 6783 5120 6828 5148
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 4356 5052 4936 5080
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 7009 5015 7067 5021
rect 7009 5012 7021 5015
rect 5868 4984 7021 5012
rect 5868 4972 5874 4984
rect 7009 4981 7021 4984
rect 7055 4981 7067 5015
rect 7009 4975 7067 4981
rect 1104 4922 21712 4944
rect 1104 4870 7851 4922
rect 7903 4870 7915 4922
rect 7967 4870 7979 4922
rect 8031 4870 8043 4922
rect 8095 4870 14720 4922
rect 14772 4870 14784 4922
rect 14836 4870 14848 4922
rect 14900 4870 14912 4922
rect 14964 4870 21712 4922
rect 1104 4848 21712 4870
rect 1489 4743 1547 4749
rect 1489 4709 1501 4743
rect 1535 4740 1547 4743
rect 2130 4740 2136 4752
rect 1535 4712 2136 4740
rect 1535 4709 1547 4712
rect 1489 4703 1547 4709
rect 2130 4700 2136 4712
rect 2188 4700 2194 4752
rect 4798 4700 4804 4752
rect 4856 4740 4862 4752
rect 4985 4743 5043 4749
rect 4985 4740 4997 4743
rect 4856 4712 4997 4740
rect 4856 4700 4862 4712
rect 4985 4709 4997 4712
rect 5031 4709 5043 4743
rect 4985 4703 5043 4709
rect 1394 4632 1400 4684
rect 1452 4672 1458 4684
rect 1946 4672 1952 4684
rect 1452 4644 1952 4672
rect 1452 4632 1458 4644
rect 1946 4632 1952 4644
rect 2004 4672 2010 4684
rect 2317 4675 2375 4681
rect 2317 4672 2329 4675
rect 2004 4644 2329 4672
rect 2004 4632 2010 4644
rect 2317 4641 2329 4644
rect 2363 4641 2375 4675
rect 2317 4635 2375 4641
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4672 2559 4675
rect 2682 4672 2688 4684
rect 2547 4644 2688 4672
rect 2547 4641 2559 4644
rect 2501 4635 2559 4641
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 4246 4632 4252 4684
rect 4304 4672 4310 4684
rect 4525 4675 4583 4681
rect 4525 4672 4537 4675
rect 4304 4644 4537 4672
rect 4304 4632 4310 4644
rect 4525 4641 4537 4644
rect 4571 4641 4583 4675
rect 5810 4672 5816 4684
rect 5771 4644 5816 4672
rect 4525 4635 4583 4641
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 5902 4632 5908 4684
rect 5960 4672 5966 4684
rect 6917 4675 6975 4681
rect 6917 4672 6929 4675
rect 5960 4644 6929 4672
rect 5960 4632 5966 4644
rect 6917 4641 6929 4644
rect 6963 4641 6975 4675
rect 6917 4635 6975 4641
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4573 2099 4607
rect 4430 4604 4436 4616
rect 4391 4576 4436 4604
rect 2041 4567 2099 4573
rect 2056 4536 2084 4567
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 3418 4536 3424 4548
rect 2056 4508 3424 4536
rect 3418 4496 3424 4508
rect 3476 4496 3482 4548
rect 5994 4468 6000 4480
rect 5955 4440 6000 4468
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 6086 4428 6092 4480
rect 6144 4468 6150 4480
rect 7101 4471 7159 4477
rect 7101 4468 7113 4471
rect 6144 4440 7113 4468
rect 6144 4428 6150 4440
rect 7101 4437 7113 4440
rect 7147 4437 7159 4471
rect 7101 4431 7159 4437
rect 1104 4378 21712 4400
rect 1104 4326 4416 4378
rect 4468 4326 4480 4378
rect 4532 4326 4544 4378
rect 4596 4326 4608 4378
rect 4660 4326 11286 4378
rect 11338 4326 11350 4378
rect 11402 4326 11414 4378
rect 11466 4326 11478 4378
rect 11530 4326 18155 4378
rect 18207 4326 18219 4378
rect 18271 4326 18283 4378
rect 18335 4326 18347 4378
rect 18399 4326 21712 4378
rect 1104 4304 21712 4326
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4060 2283 4063
rect 2314 4060 2320 4072
rect 2271 4032 2320 4060
rect 2271 4029 2283 4032
rect 2225 4023 2283 4029
rect 2314 4020 2320 4032
rect 2372 4020 2378 4072
rect 3050 4020 3056 4072
rect 3108 4060 3114 4072
rect 3329 4063 3387 4069
rect 3329 4060 3341 4063
rect 3108 4032 3341 4060
rect 3108 4020 3114 4032
rect 3329 4029 3341 4032
rect 3375 4029 3387 4063
rect 3329 4023 3387 4029
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4060 4859 4063
rect 5994 4060 6000 4072
rect 4847 4032 6000 4060
rect 4847 4029 4859 4032
rect 4801 4023 4859 4029
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 2406 3924 2412 3936
rect 2367 3896 2412 3924
rect 2406 3884 2412 3896
rect 2464 3884 2470 3936
rect 3510 3924 3516 3936
rect 3471 3896 3516 3924
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 4982 3924 4988 3936
rect 4943 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 1104 3834 21712 3856
rect 1104 3782 7851 3834
rect 7903 3782 7915 3834
rect 7967 3782 7979 3834
rect 8031 3782 8043 3834
rect 8095 3782 14720 3834
rect 14772 3782 14784 3834
rect 14836 3782 14848 3834
rect 14900 3782 14912 3834
rect 14964 3782 21712 3834
rect 1104 3760 21712 3782
rect 2409 3723 2467 3729
rect 2409 3689 2421 3723
rect 2455 3720 2467 3723
rect 2498 3720 2504 3732
rect 2455 3692 2504 3720
rect 2455 3689 2467 3692
rect 2409 3683 2467 3689
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 4706 3680 4712 3732
rect 4764 3720 4770 3732
rect 4985 3723 5043 3729
rect 4985 3720 4997 3723
rect 4764 3692 4997 3720
rect 4764 3680 4770 3692
rect 4985 3689 4997 3692
rect 5031 3689 5043 3723
rect 4985 3683 5043 3689
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3584 2283 3587
rect 3142 3584 3148 3596
rect 2271 3556 3148 3584
rect 2271 3553 2283 3556
rect 2225 3547 2283 3553
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 4801 3587 4859 3593
rect 4801 3553 4813 3587
rect 4847 3584 4859 3587
rect 6086 3584 6092 3596
rect 4847 3556 6092 3584
rect 4847 3553 4859 3556
rect 4801 3547 4859 3553
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 1104 3290 21712 3312
rect 1104 3238 4416 3290
rect 4468 3238 4480 3290
rect 4532 3238 4544 3290
rect 4596 3238 4608 3290
rect 4660 3238 11286 3290
rect 11338 3238 11350 3290
rect 11402 3238 11414 3290
rect 11466 3238 11478 3290
rect 11530 3238 18155 3290
rect 18207 3238 18219 3290
rect 18271 3238 18283 3290
rect 18335 3238 18347 3290
rect 18399 3238 21712 3290
rect 1104 3216 21712 3238
rect 2409 3179 2467 3185
rect 2409 3145 2421 3179
rect 2455 3176 2467 3179
rect 2590 3176 2596 3188
rect 2455 3148 2596 3176
rect 2455 3145 2467 3148
rect 2409 3139 2467 3145
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 3418 3176 3424 3188
rect 3379 3148 3424 3176
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 2222 2972 2228 2984
rect 2183 2944 2228 2972
rect 2222 2932 2228 2944
rect 2280 2932 2286 2984
rect 3326 2972 3332 2984
rect 3287 2944 3332 2972
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 1104 2746 21712 2768
rect 1104 2694 7851 2746
rect 7903 2694 7915 2746
rect 7967 2694 7979 2746
rect 8031 2694 8043 2746
rect 8095 2694 14720 2746
rect 14772 2694 14784 2746
rect 14836 2694 14848 2746
rect 14900 2694 14912 2746
rect 14964 2694 21712 2746
rect 1104 2672 21712 2694
rect 2038 2632 2044 2644
rect 1999 2604 2044 2632
rect 2038 2592 2044 2604
rect 2096 2592 2102 2644
rect 4062 2592 4068 2644
rect 4120 2632 4126 2644
rect 19242 2632 19248 2644
rect 4120 2604 19248 2632
rect 4120 2592 4126 2604
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 2866 2496 2872 2508
rect 1995 2468 2872 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 1104 2202 21712 2224
rect 1104 2150 4416 2202
rect 4468 2150 4480 2202
rect 4532 2150 4544 2202
rect 4596 2150 4608 2202
rect 4660 2150 11286 2202
rect 11338 2150 11350 2202
rect 11402 2150 11414 2202
rect 11466 2150 11478 2202
rect 11530 2150 18155 2202
rect 18207 2150 18219 2202
rect 18271 2150 18283 2202
rect 18335 2150 18347 2202
rect 18399 2150 21712 2202
rect 1104 2128 21712 2150
rect 20714 892 20720 944
rect 20772 932 20778 944
rect 21358 932 21364 944
rect 20772 904 21364 932
rect 20772 892 20778 904
rect 21358 892 21364 904
rect 21416 892 21422 944
<< via1 >>
rect 7851 22278 7903 22330
rect 7915 22278 7967 22330
rect 7979 22278 8031 22330
rect 8043 22278 8095 22330
rect 14720 22278 14772 22330
rect 14784 22278 14836 22330
rect 14848 22278 14900 22330
rect 14912 22278 14964 22330
rect 4416 21734 4468 21786
rect 4480 21734 4532 21786
rect 4544 21734 4596 21786
rect 4608 21734 4660 21786
rect 11286 21734 11338 21786
rect 11350 21734 11402 21786
rect 11414 21734 11466 21786
rect 11478 21734 11530 21786
rect 18155 21734 18207 21786
rect 18219 21734 18271 21786
rect 18283 21734 18335 21786
rect 18347 21734 18399 21786
rect 19248 21496 19300 21548
rect 20168 21471 20220 21480
rect 20168 21437 20177 21471
rect 20177 21437 20211 21471
rect 20211 21437 20220 21471
rect 20168 21428 20220 21437
rect 20444 21335 20496 21344
rect 20444 21301 20453 21335
rect 20453 21301 20487 21335
rect 20487 21301 20496 21335
rect 20444 21292 20496 21301
rect 7851 21190 7903 21242
rect 7915 21190 7967 21242
rect 7979 21190 8031 21242
rect 8043 21190 8095 21242
rect 14720 21190 14772 21242
rect 14784 21190 14836 21242
rect 14848 21190 14900 21242
rect 14912 21190 14964 21242
rect 19064 21131 19116 21140
rect 19064 21097 19073 21131
rect 19073 21097 19107 21131
rect 19107 21097 19116 21131
rect 19064 21088 19116 21097
rect 19248 20952 19300 21004
rect 19616 20952 19668 21004
rect 19892 20952 19944 21004
rect 21364 20952 21416 21004
rect 19524 20927 19576 20936
rect 19524 20893 19533 20927
rect 19533 20893 19567 20927
rect 19567 20893 19576 20927
rect 19524 20884 19576 20893
rect 4416 20646 4468 20698
rect 4480 20646 4532 20698
rect 4544 20646 4596 20698
rect 4608 20646 4660 20698
rect 11286 20646 11338 20698
rect 11350 20646 11402 20698
rect 11414 20646 11466 20698
rect 11478 20646 11530 20698
rect 18155 20646 18207 20698
rect 18219 20646 18271 20698
rect 18283 20646 18335 20698
rect 18347 20646 18399 20698
rect 20168 20476 20220 20528
rect 19892 20383 19944 20392
rect 19892 20349 19901 20383
rect 19901 20349 19935 20383
rect 19935 20349 19944 20383
rect 19892 20340 19944 20349
rect 19616 20272 19668 20324
rect 20720 20340 20772 20392
rect 7851 20102 7903 20154
rect 7915 20102 7967 20154
rect 7979 20102 8031 20154
rect 8043 20102 8095 20154
rect 14720 20102 14772 20154
rect 14784 20102 14836 20154
rect 14848 20102 14900 20154
rect 14912 20102 14964 20154
rect 19616 19864 19668 19916
rect 19892 19796 19944 19848
rect 19524 19660 19576 19712
rect 4416 19558 4468 19610
rect 4480 19558 4532 19610
rect 4544 19558 4596 19610
rect 4608 19558 4660 19610
rect 11286 19558 11338 19610
rect 11350 19558 11402 19610
rect 11414 19558 11466 19610
rect 11478 19558 11530 19610
rect 18155 19558 18207 19610
rect 18219 19558 18271 19610
rect 18283 19558 18335 19610
rect 18347 19558 18399 19610
rect 4252 19320 4304 19372
rect 5172 19320 5224 19372
rect 18880 19295 18932 19304
rect 18880 19261 18889 19295
rect 18889 19261 18923 19295
rect 18923 19261 18932 19295
rect 18880 19252 18932 19261
rect 18972 19295 19024 19304
rect 18972 19261 19001 19295
rect 19001 19261 19024 19295
rect 18972 19252 19024 19261
rect 19340 19184 19392 19236
rect 7851 19014 7903 19066
rect 7915 19014 7967 19066
rect 7979 19014 8031 19066
rect 8043 19014 8095 19066
rect 14720 19014 14772 19066
rect 14784 19014 14836 19066
rect 14848 19014 14900 19066
rect 14912 19014 14964 19066
rect 19248 18912 19300 18964
rect 18972 18844 19024 18896
rect 19248 18819 19300 18828
rect 19248 18785 19257 18819
rect 19257 18785 19291 18819
rect 19291 18785 19300 18819
rect 19248 18776 19300 18785
rect 19340 18751 19392 18760
rect 19340 18717 19349 18751
rect 19349 18717 19383 18751
rect 19383 18717 19392 18751
rect 19340 18708 19392 18717
rect 18880 18640 18932 18692
rect 4416 18470 4468 18522
rect 4480 18470 4532 18522
rect 4544 18470 4596 18522
rect 4608 18470 4660 18522
rect 11286 18470 11338 18522
rect 11350 18470 11402 18522
rect 11414 18470 11466 18522
rect 11478 18470 11530 18522
rect 18155 18470 18207 18522
rect 18219 18470 18271 18522
rect 18283 18470 18335 18522
rect 18347 18470 18399 18522
rect 18972 18232 19024 18284
rect 18880 18207 18932 18216
rect 18880 18173 18889 18207
rect 18889 18173 18923 18207
rect 18923 18173 18932 18207
rect 18880 18164 18932 18173
rect 19800 18071 19852 18080
rect 19800 18037 19809 18071
rect 19809 18037 19843 18071
rect 19843 18037 19852 18071
rect 19800 18028 19852 18037
rect 7851 17926 7903 17978
rect 7915 17926 7967 17978
rect 7979 17926 8031 17978
rect 8043 17926 8095 17978
rect 14720 17926 14772 17978
rect 14784 17926 14836 17978
rect 14848 17926 14900 17978
rect 14912 17926 14964 17978
rect 19892 17799 19944 17808
rect 19340 17731 19392 17740
rect 19340 17697 19349 17731
rect 19349 17697 19383 17731
rect 19383 17697 19392 17731
rect 19340 17688 19392 17697
rect 19892 17765 19901 17799
rect 19901 17765 19935 17799
rect 19935 17765 19944 17799
rect 19892 17756 19944 17765
rect 19800 17688 19852 17740
rect 4416 17382 4468 17434
rect 4480 17382 4532 17434
rect 4544 17382 4596 17434
rect 4608 17382 4660 17434
rect 11286 17382 11338 17434
rect 11350 17382 11402 17434
rect 11414 17382 11466 17434
rect 11478 17382 11530 17434
rect 18155 17382 18207 17434
rect 18219 17382 18271 17434
rect 18283 17382 18335 17434
rect 18347 17382 18399 17434
rect 19340 17280 19392 17332
rect 19248 17119 19300 17128
rect 19248 17085 19257 17119
rect 19257 17085 19291 17119
rect 19291 17085 19300 17119
rect 19248 17076 19300 17085
rect 7851 16838 7903 16890
rect 7915 16838 7967 16890
rect 7979 16838 8031 16890
rect 8043 16838 8095 16890
rect 14720 16838 14772 16890
rect 14784 16838 14836 16890
rect 14848 16838 14900 16890
rect 14912 16838 14964 16890
rect 17776 16736 17828 16788
rect 17868 16600 17920 16652
rect 4416 16294 4468 16346
rect 4480 16294 4532 16346
rect 4544 16294 4596 16346
rect 4608 16294 4660 16346
rect 11286 16294 11338 16346
rect 11350 16294 11402 16346
rect 11414 16294 11466 16346
rect 11478 16294 11530 16346
rect 18155 16294 18207 16346
rect 18219 16294 18271 16346
rect 18283 16294 18335 16346
rect 18347 16294 18399 16346
rect 19248 16192 19300 16244
rect 16212 16099 16264 16108
rect 16212 16065 16221 16099
rect 16221 16065 16255 16099
rect 16255 16065 16264 16099
rect 16212 16056 16264 16065
rect 16396 16099 16448 16108
rect 16396 16065 16405 16099
rect 16405 16065 16439 16099
rect 16439 16065 16448 16099
rect 16396 16056 16448 16065
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 16488 16031 16540 16040
rect 16488 15997 16497 16031
rect 16497 15997 16531 16031
rect 16531 15997 16540 16031
rect 16488 15988 16540 15997
rect 7851 15750 7903 15802
rect 7915 15750 7967 15802
rect 7979 15750 8031 15802
rect 8043 15750 8095 15802
rect 14720 15750 14772 15802
rect 14784 15750 14836 15802
rect 14848 15750 14900 15802
rect 14912 15750 14964 15802
rect 16396 15648 16448 15700
rect 17868 15648 17920 15700
rect 15844 15580 15896 15632
rect 15936 15512 15988 15564
rect 16396 15512 16448 15564
rect 17776 15555 17828 15564
rect 17776 15521 17785 15555
rect 17785 15521 17819 15555
rect 17819 15521 17828 15555
rect 17776 15512 17828 15521
rect 15844 15444 15896 15496
rect 16120 15308 16172 15360
rect 16948 15308 17000 15360
rect 17040 15308 17092 15360
rect 4416 15206 4468 15258
rect 4480 15206 4532 15258
rect 4544 15206 4596 15258
rect 4608 15206 4660 15258
rect 11286 15206 11338 15258
rect 11350 15206 11402 15258
rect 11414 15206 11466 15258
rect 11478 15206 11530 15258
rect 18155 15206 18207 15258
rect 18219 15206 18271 15258
rect 18283 15206 18335 15258
rect 18347 15206 18399 15258
rect 16212 15104 16264 15156
rect 15844 14943 15896 14952
rect 15844 14909 15853 14943
rect 15853 14909 15887 14943
rect 15887 14909 15896 14943
rect 15844 14900 15896 14909
rect 15936 14943 15988 14952
rect 15936 14909 15945 14943
rect 15945 14909 15979 14943
rect 15979 14909 15988 14943
rect 15936 14900 15988 14909
rect 7851 14662 7903 14714
rect 7915 14662 7967 14714
rect 7979 14662 8031 14714
rect 8043 14662 8095 14714
rect 14720 14662 14772 14714
rect 14784 14662 14836 14714
rect 14848 14662 14900 14714
rect 14912 14662 14964 14714
rect 16580 14560 16632 14612
rect 17040 14560 17092 14612
rect 18512 14492 18564 14544
rect 14556 14424 14608 14476
rect 16580 14424 16632 14476
rect 16948 14467 17000 14476
rect 16948 14433 16957 14467
rect 16957 14433 16991 14467
rect 16991 14433 17000 14467
rect 16948 14424 17000 14433
rect 17040 14467 17092 14476
rect 17040 14433 17049 14467
rect 17049 14433 17083 14467
rect 17083 14433 17092 14467
rect 17040 14424 17092 14433
rect 14372 14220 14424 14272
rect 4416 14118 4468 14170
rect 4480 14118 4532 14170
rect 4544 14118 4596 14170
rect 4608 14118 4660 14170
rect 11286 14118 11338 14170
rect 11350 14118 11402 14170
rect 11414 14118 11466 14170
rect 11478 14118 11530 14170
rect 18155 14118 18207 14170
rect 18219 14118 18271 14170
rect 18283 14118 18335 14170
rect 18347 14118 18399 14170
rect 14556 14059 14608 14068
rect 14556 14025 14565 14059
rect 14565 14025 14599 14059
rect 14599 14025 14608 14059
rect 14556 14016 14608 14025
rect 12440 13880 12492 13932
rect 13452 13812 13504 13864
rect 13636 13812 13688 13864
rect 13360 13744 13412 13796
rect 13728 13676 13780 13728
rect 7851 13574 7903 13626
rect 7915 13574 7967 13626
rect 7979 13574 8031 13626
rect 8043 13574 8095 13626
rect 14720 13574 14772 13626
rect 14784 13574 14836 13626
rect 14848 13574 14900 13626
rect 14912 13574 14964 13626
rect 16120 13472 16172 13524
rect 13268 13379 13320 13388
rect 13268 13345 13277 13379
rect 13277 13345 13311 13379
rect 13311 13345 13320 13379
rect 13268 13336 13320 13345
rect 13452 13336 13504 13388
rect 13728 13379 13780 13388
rect 13728 13345 13737 13379
rect 13737 13345 13771 13379
rect 13771 13345 13780 13379
rect 13728 13336 13780 13345
rect 13360 13311 13412 13320
rect 13360 13277 13369 13311
rect 13369 13277 13403 13311
rect 13403 13277 13412 13311
rect 13360 13268 13412 13277
rect 4416 13030 4468 13082
rect 4480 13030 4532 13082
rect 4544 13030 4596 13082
rect 4608 13030 4660 13082
rect 11286 13030 11338 13082
rect 11350 13030 11402 13082
rect 11414 13030 11466 13082
rect 11478 13030 11530 13082
rect 18155 13030 18207 13082
rect 18219 13030 18271 13082
rect 18283 13030 18335 13082
rect 18347 13030 18399 13082
rect 13544 12724 13596 12776
rect 14004 12724 14056 12776
rect 14372 12724 14424 12776
rect 19156 12656 19208 12708
rect 13820 12588 13872 12640
rect 7851 12486 7903 12538
rect 7915 12486 7967 12538
rect 7979 12486 8031 12538
rect 8043 12486 8095 12538
rect 14720 12486 14772 12538
rect 14784 12486 14836 12538
rect 14848 12486 14900 12538
rect 14912 12486 14964 12538
rect 13452 12291 13504 12300
rect 13452 12257 13461 12291
rect 13461 12257 13495 12291
rect 13495 12257 13504 12291
rect 13452 12248 13504 12257
rect 13728 12316 13780 12368
rect 14004 12359 14056 12368
rect 14004 12325 14013 12359
rect 14013 12325 14047 12359
rect 14047 12325 14056 12359
rect 14004 12316 14056 12325
rect 12716 12223 12768 12232
rect 12716 12189 12725 12223
rect 12725 12189 12759 12223
rect 12759 12189 12768 12223
rect 12716 12180 12768 12189
rect 4416 11942 4468 11994
rect 4480 11942 4532 11994
rect 4544 11942 4596 11994
rect 4608 11942 4660 11994
rect 11286 11942 11338 11994
rect 11350 11942 11402 11994
rect 11414 11942 11466 11994
rect 11478 11942 11530 11994
rect 18155 11942 18207 11994
rect 18219 11942 18271 11994
rect 18283 11942 18335 11994
rect 18347 11942 18399 11994
rect 13544 11883 13596 11892
rect 13544 11849 13553 11883
rect 13553 11849 13587 11883
rect 13587 11849 13596 11883
rect 13544 11840 13596 11849
rect 10508 11679 10560 11688
rect 10508 11645 10517 11679
rect 10517 11645 10551 11679
rect 10551 11645 10560 11679
rect 10508 11636 10560 11645
rect 13820 11636 13872 11688
rect 11704 11500 11756 11552
rect 7851 11398 7903 11450
rect 7915 11398 7967 11450
rect 7979 11398 8031 11450
rect 8043 11398 8095 11450
rect 14720 11398 14772 11450
rect 14784 11398 14836 11450
rect 14848 11398 14900 11450
rect 14912 11398 14964 11450
rect 10600 11296 10652 11348
rect 13636 11296 13688 11348
rect 11152 11160 11204 11212
rect 13360 11203 13412 11212
rect 10416 11092 10468 11144
rect 13360 11169 13369 11203
rect 13369 11169 13403 11203
rect 13403 11169 13412 11203
rect 13360 11160 13412 11169
rect 9680 11024 9732 11076
rect 4416 10854 4468 10906
rect 4480 10854 4532 10906
rect 4544 10854 4596 10906
rect 4608 10854 4660 10906
rect 11286 10854 11338 10906
rect 11350 10854 11402 10906
rect 11414 10854 11466 10906
rect 11478 10854 11530 10906
rect 18155 10854 18207 10906
rect 18219 10854 18271 10906
rect 18283 10854 18335 10906
rect 18347 10854 18399 10906
rect 10508 10752 10560 10804
rect 9680 10548 9732 10600
rect 9956 10548 10008 10600
rect 10232 10591 10284 10600
rect 10232 10557 10241 10591
rect 10241 10557 10275 10591
rect 10275 10557 10284 10591
rect 10232 10548 10284 10557
rect 10508 10480 10560 10532
rect 7851 10310 7903 10362
rect 7915 10310 7967 10362
rect 7979 10310 8031 10362
rect 8043 10310 8095 10362
rect 14720 10310 14772 10362
rect 14784 10310 14836 10362
rect 14848 10310 14900 10362
rect 14912 10310 14964 10362
rect 11152 10208 11204 10260
rect 10692 10072 10744 10124
rect 11152 10072 11204 10124
rect 11704 10072 11756 10124
rect 19248 10004 19300 10056
rect 4416 9766 4468 9818
rect 4480 9766 4532 9818
rect 4544 9766 4596 9818
rect 4608 9766 4660 9818
rect 11286 9766 11338 9818
rect 11350 9766 11402 9818
rect 11414 9766 11466 9818
rect 11478 9766 11530 9818
rect 18155 9766 18207 9818
rect 18219 9766 18271 9818
rect 18283 9766 18335 9818
rect 18347 9766 18399 9818
rect 11152 9664 11204 9716
rect 5172 9596 5224 9648
rect 5356 9596 5408 9648
rect 9956 9571 10008 9580
rect 9956 9537 9965 9571
rect 9965 9537 9999 9571
rect 9999 9537 10008 9571
rect 9956 9528 10008 9537
rect 10140 9460 10192 9512
rect 10784 9392 10836 9444
rect 7851 9222 7903 9274
rect 7915 9222 7967 9274
rect 7979 9222 8031 9274
rect 8043 9222 8095 9274
rect 14720 9222 14772 9274
rect 14784 9222 14836 9274
rect 14848 9222 14900 9274
rect 14912 9222 14964 9274
rect 13360 9120 13412 9172
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 10416 9027 10468 9036
rect 10416 8993 10425 9027
rect 10425 8993 10459 9027
rect 10459 8993 10468 9027
rect 10416 8984 10468 8993
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 9956 8848 10008 8900
rect 9588 8780 9640 8832
rect 4416 8678 4468 8730
rect 4480 8678 4532 8730
rect 4544 8678 4596 8730
rect 4608 8678 4660 8730
rect 11286 8678 11338 8730
rect 11350 8678 11402 8730
rect 11414 8678 11466 8730
rect 11478 8678 11530 8730
rect 18155 8678 18207 8730
rect 18219 8678 18271 8730
rect 18283 8678 18335 8730
rect 18347 8678 18399 8730
rect 5908 8576 5960 8628
rect 10692 8619 10744 8628
rect 10692 8585 10701 8619
rect 10701 8585 10735 8619
rect 10735 8585 10744 8619
rect 10692 8576 10744 8585
rect 3056 8508 3108 8560
rect 6920 8508 6972 8560
rect 2596 8372 2648 8424
rect 8668 8372 8720 8424
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8760 8372 8812 8381
rect 10600 8372 10652 8424
rect 7851 8134 7903 8186
rect 7915 8134 7967 8186
rect 7979 8134 8031 8186
rect 8043 8134 8095 8186
rect 14720 8134 14772 8186
rect 14784 8134 14836 8186
rect 14848 8134 14900 8186
rect 14912 8134 14964 8186
rect 7656 8032 7708 8084
rect 2504 7896 2556 7948
rect 4712 7896 4764 7948
rect 6920 7896 6972 7948
rect 7104 7896 7156 7948
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 2320 7692 2372 7744
rect 6828 7692 6880 7744
rect 7472 7692 7524 7744
rect 4416 7590 4468 7642
rect 4480 7590 4532 7642
rect 4544 7590 4596 7642
rect 4608 7590 4660 7642
rect 11286 7590 11338 7642
rect 11350 7590 11402 7642
rect 11414 7590 11466 7642
rect 11478 7590 11530 7642
rect 18155 7590 18207 7642
rect 18219 7590 18271 7642
rect 18283 7590 18335 7642
rect 18347 7590 18399 7642
rect 8668 7488 8720 7540
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 2412 7284 2464 7336
rect 3516 7284 3568 7336
rect 4988 7284 5040 7336
rect 8208 7284 8260 7336
rect 2228 7148 2280 7200
rect 3148 7148 3200 7200
rect 4804 7148 4856 7200
rect 7748 7148 7800 7200
rect 9588 7284 9640 7336
rect 8852 7191 8904 7200
rect 8852 7157 8861 7191
rect 8861 7157 8895 7191
rect 8895 7157 8904 7191
rect 8852 7148 8904 7157
rect 7851 7046 7903 7098
rect 7915 7046 7967 7098
rect 7979 7046 8031 7098
rect 8043 7046 8095 7098
rect 14720 7046 14772 7098
rect 14784 7046 14836 7098
rect 14848 7046 14900 7098
rect 14912 7046 14964 7098
rect 8208 6987 8260 6996
rect 8208 6953 8217 6987
rect 8217 6953 8251 6987
rect 8251 6953 8260 6987
rect 8208 6944 8260 6953
rect 8852 6944 8904 6996
rect 18052 6944 18104 6996
rect 7288 6876 7340 6928
rect 7840 6876 7892 6928
rect 2228 6851 2280 6860
rect 2228 6817 2237 6851
rect 2237 6817 2271 6851
rect 2271 6817 2280 6851
rect 2228 6808 2280 6817
rect 4804 6851 4856 6860
rect 4804 6817 4813 6851
rect 4813 6817 4847 6851
rect 4847 6817 4856 6851
rect 4804 6808 4856 6817
rect 5908 6851 5960 6860
rect 5908 6817 5917 6851
rect 5917 6817 5951 6851
rect 5951 6817 5960 6851
rect 5908 6808 5960 6817
rect 7104 6808 7156 6860
rect 7288 6740 7340 6792
rect 3332 6604 3384 6656
rect 4896 6604 4948 6656
rect 7656 6604 7708 6656
rect 4416 6502 4468 6554
rect 4480 6502 4532 6554
rect 4544 6502 4596 6554
rect 4608 6502 4660 6554
rect 11286 6502 11338 6554
rect 11350 6502 11402 6554
rect 11414 6502 11466 6554
rect 11478 6502 11530 6554
rect 18155 6502 18207 6554
rect 18219 6502 18271 6554
rect 18283 6502 18335 6554
rect 18347 6502 18399 6554
rect 10416 6400 10468 6452
rect 4252 6332 4304 6384
rect 2136 6264 2188 6316
rect 2688 6264 2740 6316
rect 4804 6307 4856 6316
rect 4804 6273 4813 6307
rect 4813 6273 4847 6307
rect 4847 6273 4856 6307
rect 4804 6264 4856 6273
rect 1952 6196 2004 6248
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 2228 6128 2280 6180
rect 5356 6196 5408 6248
rect 8760 6332 8812 6384
rect 7840 6307 7892 6316
rect 7840 6273 7849 6307
rect 7849 6273 7883 6307
rect 7883 6273 7892 6307
rect 7840 6264 7892 6273
rect 5908 6128 5960 6180
rect 7104 6128 7156 6180
rect 7851 5958 7903 6010
rect 7915 5958 7967 6010
rect 7979 5958 8031 6010
rect 8043 5958 8095 6010
rect 14720 5958 14772 6010
rect 14784 5958 14836 6010
rect 14848 5958 14900 6010
rect 14912 5958 14964 6010
rect 7748 5856 7800 5908
rect 2228 5720 2280 5772
rect 1952 5652 2004 5704
rect 2688 5720 2740 5772
rect 4896 5720 4948 5772
rect 5356 5720 5408 5772
rect 7656 5763 7708 5772
rect 7656 5729 7665 5763
rect 7665 5729 7699 5763
rect 7699 5729 7708 5763
rect 7656 5720 7708 5729
rect 2872 5584 2924 5636
rect 18788 5584 18840 5636
rect 5908 5516 5960 5568
rect 4416 5414 4468 5466
rect 4480 5414 4532 5466
rect 4544 5414 4596 5466
rect 4608 5414 4660 5466
rect 11286 5414 11338 5466
rect 11350 5414 11402 5466
rect 11414 5414 11466 5466
rect 11478 5414 11530 5466
rect 18155 5414 18207 5466
rect 18219 5414 18271 5466
rect 18283 5414 18335 5466
rect 18347 5414 18399 5466
rect 5356 5355 5408 5364
rect 5356 5321 5365 5355
rect 5365 5321 5399 5355
rect 5399 5321 5408 5355
rect 5356 5312 5408 5321
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 2136 5151 2188 5160
rect 2136 5117 2145 5151
rect 2145 5117 2179 5151
rect 2179 5117 2188 5151
rect 2136 5108 2188 5117
rect 4252 5108 4304 5160
rect 4068 5040 4120 5092
rect 4436 5151 4488 5160
rect 4436 5117 4445 5151
rect 4445 5117 4479 5151
rect 4479 5117 4488 5151
rect 5264 5244 5316 5296
rect 4436 5108 4488 5117
rect 5264 5108 5316 5160
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 5816 4972 5868 5024
rect 7851 4870 7903 4922
rect 7915 4870 7967 4922
rect 7979 4870 8031 4922
rect 8043 4870 8095 4922
rect 14720 4870 14772 4922
rect 14784 4870 14836 4922
rect 14848 4870 14900 4922
rect 14912 4870 14964 4922
rect 2136 4700 2188 4752
rect 4804 4700 4856 4752
rect 1400 4632 1452 4684
rect 1952 4632 2004 4684
rect 2688 4632 2740 4684
rect 4252 4632 4304 4684
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 5908 4632 5960 4684
rect 4436 4607 4488 4616
rect 4436 4573 4445 4607
rect 4445 4573 4479 4607
rect 4479 4573 4488 4607
rect 4436 4564 4488 4573
rect 3424 4496 3476 4548
rect 6000 4471 6052 4480
rect 6000 4437 6009 4471
rect 6009 4437 6043 4471
rect 6043 4437 6052 4471
rect 6000 4428 6052 4437
rect 6092 4428 6144 4480
rect 4416 4326 4468 4378
rect 4480 4326 4532 4378
rect 4544 4326 4596 4378
rect 4608 4326 4660 4378
rect 11286 4326 11338 4378
rect 11350 4326 11402 4378
rect 11414 4326 11466 4378
rect 11478 4326 11530 4378
rect 18155 4326 18207 4378
rect 18219 4326 18271 4378
rect 18283 4326 18335 4378
rect 18347 4326 18399 4378
rect 2320 4020 2372 4072
rect 3056 4020 3108 4072
rect 6000 4020 6052 4072
rect 2412 3927 2464 3936
rect 2412 3893 2421 3927
rect 2421 3893 2455 3927
rect 2455 3893 2464 3927
rect 2412 3884 2464 3893
rect 3516 3927 3568 3936
rect 3516 3893 3525 3927
rect 3525 3893 3559 3927
rect 3559 3893 3568 3927
rect 3516 3884 3568 3893
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 7851 3782 7903 3834
rect 7915 3782 7967 3834
rect 7979 3782 8031 3834
rect 8043 3782 8095 3834
rect 14720 3782 14772 3834
rect 14784 3782 14836 3834
rect 14848 3782 14900 3834
rect 14912 3782 14964 3834
rect 2504 3680 2556 3732
rect 4712 3680 4764 3732
rect 3148 3544 3200 3596
rect 6092 3544 6144 3596
rect 4416 3238 4468 3290
rect 4480 3238 4532 3290
rect 4544 3238 4596 3290
rect 4608 3238 4660 3290
rect 11286 3238 11338 3290
rect 11350 3238 11402 3290
rect 11414 3238 11466 3290
rect 11478 3238 11530 3290
rect 18155 3238 18207 3290
rect 18219 3238 18271 3290
rect 18283 3238 18335 3290
rect 18347 3238 18399 3290
rect 2596 3136 2648 3188
rect 3424 3179 3476 3188
rect 3424 3145 3433 3179
rect 3433 3145 3467 3179
rect 3467 3145 3476 3179
rect 3424 3136 3476 3145
rect 2228 2975 2280 2984
rect 2228 2941 2237 2975
rect 2237 2941 2271 2975
rect 2271 2941 2280 2975
rect 2228 2932 2280 2941
rect 3332 2975 3384 2984
rect 3332 2941 3341 2975
rect 3341 2941 3375 2975
rect 3375 2941 3384 2975
rect 3332 2932 3384 2941
rect 7851 2694 7903 2746
rect 7915 2694 7967 2746
rect 7979 2694 8031 2746
rect 8043 2694 8095 2746
rect 14720 2694 14772 2746
rect 14784 2694 14836 2746
rect 14848 2694 14900 2746
rect 14912 2694 14964 2746
rect 2044 2635 2096 2644
rect 2044 2601 2053 2635
rect 2053 2601 2087 2635
rect 2087 2601 2096 2635
rect 2044 2592 2096 2601
rect 4068 2592 4120 2644
rect 19248 2592 19300 2644
rect 2872 2456 2924 2508
rect 4416 2150 4468 2202
rect 4480 2150 4532 2202
rect 4544 2150 4596 2202
rect 4608 2150 4660 2202
rect 11286 2150 11338 2202
rect 11350 2150 11402 2202
rect 11414 2150 11466 2202
rect 11478 2150 11530 2202
rect 18155 2150 18207 2202
rect 18219 2150 18271 2202
rect 18283 2150 18335 2202
rect 18347 2150 18399 2202
rect 20720 892 20772 944
rect 21364 892 21416 944
<< metal2 >>
rect 1398 24202 1454 25002
rect 4250 24202 4306 25002
rect 7102 24202 7158 25002
rect 9954 24202 10010 25002
rect 12806 24202 12862 25002
rect 15658 24202 15714 25002
rect 18510 24202 18566 25002
rect 21362 24202 21418 25002
rect 1412 24154 1440 24202
rect 1412 24126 2360 24154
rect 2332 9602 2360 24126
rect 4264 19378 4292 24202
rect 7116 24154 7144 24202
rect 9968 24154 9996 24202
rect 12820 24154 12848 24202
rect 7116 24126 7328 24154
rect 9968 24126 10272 24154
rect 4390 21788 4686 21808
rect 4446 21786 4470 21788
rect 4526 21786 4550 21788
rect 4606 21786 4630 21788
rect 4468 21734 4470 21786
rect 4532 21734 4544 21786
rect 4606 21734 4608 21786
rect 4446 21732 4470 21734
rect 4526 21732 4550 21734
rect 4606 21732 4630 21734
rect 4390 21712 4686 21732
rect 4390 20700 4686 20720
rect 4446 20698 4470 20700
rect 4526 20698 4550 20700
rect 4606 20698 4630 20700
rect 4468 20646 4470 20698
rect 4532 20646 4544 20698
rect 4606 20646 4608 20698
rect 4446 20644 4470 20646
rect 4526 20644 4550 20646
rect 4606 20644 4630 20646
rect 4390 20624 4686 20644
rect 4390 19612 4686 19632
rect 4446 19610 4470 19612
rect 4526 19610 4550 19612
rect 4606 19610 4630 19612
rect 4468 19558 4470 19610
rect 4532 19558 4544 19610
rect 4606 19558 4608 19610
rect 4446 19556 4470 19558
rect 4526 19556 4550 19558
rect 4606 19556 4630 19558
rect 4390 19536 4686 19556
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 4390 18524 4686 18544
rect 4446 18522 4470 18524
rect 4526 18522 4550 18524
rect 4606 18522 4630 18524
rect 4468 18470 4470 18522
rect 4532 18470 4544 18522
rect 4606 18470 4608 18522
rect 4446 18468 4470 18470
rect 4526 18468 4550 18470
rect 4606 18468 4630 18470
rect 4390 18448 4686 18468
rect 4390 17436 4686 17456
rect 4446 17434 4470 17436
rect 4526 17434 4550 17436
rect 4606 17434 4630 17436
rect 4468 17382 4470 17434
rect 4532 17382 4544 17434
rect 4606 17382 4608 17434
rect 4446 17380 4470 17382
rect 4526 17380 4550 17382
rect 4606 17380 4630 17382
rect 4390 17360 4686 17380
rect 4390 16348 4686 16368
rect 4446 16346 4470 16348
rect 4526 16346 4550 16348
rect 4606 16346 4630 16348
rect 4468 16294 4470 16346
rect 4532 16294 4544 16346
rect 4606 16294 4608 16346
rect 4446 16292 4470 16294
rect 4526 16292 4550 16294
rect 4606 16292 4630 16294
rect 4390 16272 4686 16292
rect 4390 15260 4686 15280
rect 4446 15258 4470 15260
rect 4526 15258 4550 15260
rect 4606 15258 4630 15260
rect 4468 15206 4470 15258
rect 4532 15206 4544 15258
rect 4606 15206 4608 15258
rect 4446 15204 4470 15206
rect 4526 15204 4550 15206
rect 4606 15204 4630 15206
rect 4390 15184 4686 15204
rect 4390 14172 4686 14192
rect 4446 14170 4470 14172
rect 4526 14170 4550 14172
rect 4606 14170 4630 14172
rect 4468 14118 4470 14170
rect 4532 14118 4544 14170
rect 4606 14118 4608 14170
rect 4446 14116 4470 14118
rect 4526 14116 4550 14118
rect 4606 14116 4630 14118
rect 4390 14096 4686 14116
rect 4390 13084 4686 13104
rect 4446 13082 4470 13084
rect 4526 13082 4550 13084
rect 4606 13082 4630 13084
rect 4468 13030 4470 13082
rect 4532 13030 4544 13082
rect 4606 13030 4608 13082
rect 4446 13028 4470 13030
rect 4526 13028 4550 13030
rect 4606 13028 4630 13030
rect 4390 13008 4686 13028
rect 2870 12608 2926 12617
rect 2870 12543 2926 12552
rect 2148 9574 2360 9602
rect 2148 6322 2176 9574
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2240 6866 2268 7142
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1964 5710 1992 6190
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 2240 5778 2268 6122
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1964 4690 1992 5646
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1412 800 1440 4626
rect 2056 2650 2084 5170
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 2148 4758 2176 5102
rect 2136 4752 2188 4758
rect 2136 4694 2188 4700
rect 2240 2990 2268 5714
rect 2332 4078 2360 7686
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 2424 3942 2452 7278
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2516 3738 2544 7890
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2608 3194 2636 8366
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2700 5778 2728 6258
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2700 4690 2728 5714
rect 2884 5642 2912 12543
rect 4390 11996 4686 12016
rect 4446 11994 4470 11996
rect 4526 11994 4550 11996
rect 4606 11994 4630 11996
rect 4468 11942 4470 11994
rect 4532 11942 4544 11994
rect 4606 11942 4608 11994
rect 4446 11940 4470 11942
rect 4526 11940 4550 11942
rect 4606 11940 4630 11942
rect 4390 11920 4686 11940
rect 4390 10908 4686 10928
rect 4446 10906 4470 10908
rect 4526 10906 4550 10908
rect 4606 10906 4630 10908
rect 4468 10854 4470 10906
rect 4532 10854 4544 10906
rect 4606 10854 4608 10906
rect 4446 10852 4470 10854
rect 4526 10852 4550 10854
rect 4606 10852 4630 10854
rect 4390 10832 4686 10852
rect 4390 9820 4686 9840
rect 4446 9818 4470 9820
rect 4526 9818 4550 9820
rect 4606 9818 4630 9820
rect 4468 9766 4470 9818
rect 4532 9766 4544 9818
rect 4606 9766 4608 9818
rect 4446 9764 4470 9766
rect 4526 9764 4550 9766
rect 4606 9764 4630 9766
rect 4390 9744 4686 9764
rect 5184 9654 5212 19314
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 4390 8732 4686 8752
rect 4446 8730 4470 8732
rect 4526 8730 4550 8732
rect 4606 8730 4630 8732
rect 4468 8678 4470 8730
rect 4532 8678 4544 8730
rect 4606 8678 4608 8730
rect 4446 8676 4470 8678
rect 4526 8676 4550 8678
rect 4606 8676 4630 8678
rect 4390 8656 4686 8676
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 2884 2514 2912 5578
rect 3068 4078 3096 8502
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4390 7644 4686 7664
rect 4446 7642 4470 7644
rect 4526 7642 4550 7644
rect 4606 7642 4630 7644
rect 4468 7590 4470 7642
rect 4532 7590 4544 7642
rect 4606 7590 4608 7642
rect 4446 7588 4470 7590
rect 4526 7588 4550 7590
rect 4606 7588 4630 7590
rect 4390 7568 4686 7588
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 3160 3602 3188 7142
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3344 2990 3372 6598
rect 3424 4548 3476 4554
rect 3424 4490 3476 4496
rect 3436 3194 3464 4490
rect 3528 3942 3556 7278
rect 4390 6556 4686 6576
rect 4446 6554 4470 6556
rect 4526 6554 4550 6556
rect 4606 6554 4630 6556
rect 4468 6502 4470 6554
rect 4532 6502 4544 6554
rect 4606 6502 4608 6554
rect 4446 6500 4470 6502
rect 4526 6500 4550 6502
rect 4606 6500 4630 6502
rect 4390 6480 4686 6500
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 4264 5166 4292 6326
rect 4390 5468 4686 5488
rect 4446 5466 4470 5468
rect 4526 5466 4550 5468
rect 4606 5466 4630 5468
rect 4468 5414 4470 5466
rect 4532 5414 4544 5466
rect 4606 5414 4608 5466
rect 4446 5412 4470 5414
rect 4526 5412 4550 5414
rect 4606 5412 4630 5414
rect 4390 5392 4686 5412
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 4080 2650 4108 5034
rect 4264 4690 4292 5102
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 4264 800 4292 4626
rect 4448 4622 4476 5102
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4390 4380 4686 4400
rect 4446 4378 4470 4380
rect 4526 4378 4550 4380
rect 4606 4378 4630 4380
rect 4468 4326 4470 4378
rect 4532 4326 4544 4378
rect 4606 4326 4608 4378
rect 4446 4324 4470 4326
rect 4526 4324 4550 4326
rect 4606 4324 4630 4326
rect 4390 4304 4686 4324
rect 4724 3738 4752 7890
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4816 6866 4844 7142
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 4816 4758 4844 6258
rect 4908 5778 4936 6598
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 5000 3942 5028 7278
rect 5368 6254 5396 9590
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5920 6866 5948 8570
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6932 7954 6960 8502
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5356 6248 5408 6254
rect 5276 6208 5356 6236
rect 5276 5302 5304 6208
rect 5356 6190 5408 6196
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5368 5370 5396 5714
rect 5920 5574 5948 6122
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 5276 5166 5304 5238
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5828 4690 5856 4966
rect 5920 4690 5948 5510
rect 6840 5166 6868 7686
rect 7116 6866 7144 7890
rect 7300 7886 7328 24126
rect 7825 22332 8121 22352
rect 7881 22330 7905 22332
rect 7961 22330 7985 22332
rect 8041 22330 8065 22332
rect 7903 22278 7905 22330
rect 7967 22278 7979 22330
rect 8041 22278 8043 22330
rect 7881 22276 7905 22278
rect 7961 22276 7985 22278
rect 8041 22276 8065 22278
rect 7825 22256 8121 22276
rect 7825 21244 8121 21264
rect 7881 21242 7905 21244
rect 7961 21242 7985 21244
rect 8041 21242 8065 21244
rect 7903 21190 7905 21242
rect 7967 21190 7979 21242
rect 8041 21190 8043 21242
rect 7881 21188 7905 21190
rect 7961 21188 7985 21190
rect 8041 21188 8065 21190
rect 7825 21168 8121 21188
rect 7825 20156 8121 20176
rect 7881 20154 7905 20156
rect 7961 20154 7985 20156
rect 8041 20154 8065 20156
rect 7903 20102 7905 20154
rect 7967 20102 7979 20154
rect 8041 20102 8043 20154
rect 7881 20100 7905 20102
rect 7961 20100 7985 20102
rect 8041 20100 8065 20102
rect 7825 20080 8121 20100
rect 7825 19068 8121 19088
rect 7881 19066 7905 19068
rect 7961 19066 7985 19068
rect 8041 19066 8065 19068
rect 7903 19014 7905 19066
rect 7967 19014 7979 19066
rect 8041 19014 8043 19066
rect 7881 19012 7905 19014
rect 7961 19012 7985 19014
rect 8041 19012 8065 19014
rect 7825 18992 8121 19012
rect 7825 17980 8121 18000
rect 7881 17978 7905 17980
rect 7961 17978 7985 17980
rect 8041 17978 8065 17980
rect 7903 17926 7905 17978
rect 7967 17926 7979 17978
rect 8041 17926 8043 17978
rect 7881 17924 7905 17926
rect 7961 17924 7985 17926
rect 8041 17924 8065 17926
rect 7825 17904 8121 17924
rect 7825 16892 8121 16912
rect 7881 16890 7905 16892
rect 7961 16890 7985 16892
rect 8041 16890 8065 16892
rect 7903 16838 7905 16890
rect 7967 16838 7979 16890
rect 8041 16838 8043 16890
rect 7881 16836 7905 16838
rect 7961 16836 7985 16838
rect 8041 16836 8065 16838
rect 7825 16816 8121 16836
rect 7825 15804 8121 15824
rect 7881 15802 7905 15804
rect 7961 15802 7985 15804
rect 8041 15802 8065 15804
rect 7903 15750 7905 15802
rect 7967 15750 7979 15802
rect 8041 15750 8043 15802
rect 7881 15748 7905 15750
rect 7961 15748 7985 15750
rect 8041 15748 8065 15750
rect 7825 15728 8121 15748
rect 7825 14716 8121 14736
rect 7881 14714 7905 14716
rect 7961 14714 7985 14716
rect 8041 14714 8065 14716
rect 7903 14662 7905 14714
rect 7967 14662 7979 14714
rect 8041 14662 8043 14714
rect 7881 14660 7905 14662
rect 7961 14660 7985 14662
rect 8041 14660 8065 14662
rect 7825 14640 8121 14660
rect 7825 13628 8121 13648
rect 7881 13626 7905 13628
rect 7961 13626 7985 13628
rect 8041 13626 8065 13628
rect 7903 13574 7905 13626
rect 7967 13574 7979 13626
rect 8041 13574 8043 13626
rect 7881 13572 7905 13574
rect 7961 13572 7985 13574
rect 8041 13572 8065 13574
rect 7825 13552 8121 13572
rect 7825 12540 8121 12560
rect 7881 12538 7905 12540
rect 7961 12538 7985 12540
rect 8041 12538 8065 12540
rect 7903 12486 7905 12538
rect 7967 12486 7979 12538
rect 8041 12486 8043 12538
rect 7881 12484 7905 12486
rect 7961 12484 7985 12486
rect 8041 12484 8065 12486
rect 7825 12464 8121 12484
rect 7825 11452 8121 11472
rect 7881 11450 7905 11452
rect 7961 11450 7985 11452
rect 8041 11450 8065 11452
rect 7903 11398 7905 11450
rect 7967 11398 7979 11450
rect 8041 11398 8043 11450
rect 7881 11396 7905 11398
rect 7961 11396 7985 11398
rect 8041 11396 8065 11398
rect 7825 11376 8121 11396
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 10606 9720 11018
rect 10244 10606 10272 24126
rect 12452 24126 12848 24154
rect 15672 24154 15700 24202
rect 15672 24126 16528 24154
rect 11260 21788 11556 21808
rect 11316 21786 11340 21788
rect 11396 21786 11420 21788
rect 11476 21786 11500 21788
rect 11338 21734 11340 21786
rect 11402 21734 11414 21786
rect 11476 21734 11478 21786
rect 11316 21732 11340 21734
rect 11396 21732 11420 21734
rect 11476 21732 11500 21734
rect 11260 21712 11556 21732
rect 11260 20700 11556 20720
rect 11316 20698 11340 20700
rect 11396 20698 11420 20700
rect 11476 20698 11500 20700
rect 11338 20646 11340 20698
rect 11402 20646 11414 20698
rect 11476 20646 11478 20698
rect 11316 20644 11340 20646
rect 11396 20644 11420 20646
rect 11476 20644 11500 20646
rect 11260 20624 11556 20644
rect 11260 19612 11556 19632
rect 11316 19610 11340 19612
rect 11396 19610 11420 19612
rect 11476 19610 11500 19612
rect 11338 19558 11340 19610
rect 11402 19558 11414 19610
rect 11476 19558 11478 19610
rect 11316 19556 11340 19558
rect 11396 19556 11420 19558
rect 11476 19556 11500 19558
rect 11260 19536 11556 19556
rect 11260 18524 11556 18544
rect 11316 18522 11340 18524
rect 11396 18522 11420 18524
rect 11476 18522 11500 18524
rect 11338 18470 11340 18522
rect 11402 18470 11414 18522
rect 11476 18470 11478 18522
rect 11316 18468 11340 18470
rect 11396 18468 11420 18470
rect 11476 18468 11500 18470
rect 11260 18448 11556 18468
rect 11260 17436 11556 17456
rect 11316 17434 11340 17436
rect 11396 17434 11420 17436
rect 11476 17434 11500 17436
rect 11338 17382 11340 17434
rect 11402 17382 11414 17434
rect 11476 17382 11478 17434
rect 11316 17380 11340 17382
rect 11396 17380 11420 17382
rect 11476 17380 11500 17382
rect 11260 17360 11556 17380
rect 11260 16348 11556 16368
rect 11316 16346 11340 16348
rect 11396 16346 11420 16348
rect 11476 16346 11500 16348
rect 11338 16294 11340 16346
rect 11402 16294 11414 16346
rect 11476 16294 11478 16346
rect 11316 16292 11340 16294
rect 11396 16292 11420 16294
rect 11476 16292 11500 16294
rect 11260 16272 11556 16292
rect 11260 15260 11556 15280
rect 11316 15258 11340 15260
rect 11396 15258 11420 15260
rect 11476 15258 11500 15260
rect 11338 15206 11340 15258
rect 11402 15206 11414 15258
rect 11476 15206 11478 15258
rect 11316 15204 11340 15206
rect 11396 15204 11420 15206
rect 11476 15204 11500 15206
rect 11260 15184 11556 15204
rect 11260 14172 11556 14192
rect 11316 14170 11340 14172
rect 11396 14170 11420 14172
rect 11476 14170 11500 14172
rect 11338 14118 11340 14170
rect 11402 14118 11414 14170
rect 11476 14118 11478 14170
rect 11316 14116 11340 14118
rect 11396 14116 11420 14118
rect 11476 14116 11500 14118
rect 11260 14096 11556 14116
rect 12452 13938 12480 24126
rect 14694 22332 14990 22352
rect 14750 22330 14774 22332
rect 14830 22330 14854 22332
rect 14910 22330 14934 22332
rect 14772 22278 14774 22330
rect 14836 22278 14848 22330
rect 14910 22278 14912 22330
rect 14750 22276 14774 22278
rect 14830 22276 14854 22278
rect 14910 22276 14934 22278
rect 14694 22256 14990 22276
rect 14694 21244 14990 21264
rect 14750 21242 14774 21244
rect 14830 21242 14854 21244
rect 14910 21242 14934 21244
rect 14772 21190 14774 21242
rect 14836 21190 14848 21242
rect 14910 21190 14912 21242
rect 14750 21188 14774 21190
rect 14830 21188 14854 21190
rect 14910 21188 14934 21190
rect 14694 21168 14990 21188
rect 14694 20156 14990 20176
rect 14750 20154 14774 20156
rect 14830 20154 14854 20156
rect 14910 20154 14934 20156
rect 14772 20102 14774 20154
rect 14836 20102 14848 20154
rect 14910 20102 14912 20154
rect 14750 20100 14774 20102
rect 14830 20100 14854 20102
rect 14910 20100 14934 20102
rect 14694 20080 14990 20100
rect 14694 19068 14990 19088
rect 14750 19066 14774 19068
rect 14830 19066 14854 19068
rect 14910 19066 14934 19068
rect 14772 19014 14774 19066
rect 14836 19014 14848 19066
rect 14910 19014 14912 19066
rect 14750 19012 14774 19014
rect 14830 19012 14854 19014
rect 14910 19012 14934 19014
rect 14694 18992 14990 19012
rect 14694 17980 14990 18000
rect 14750 17978 14774 17980
rect 14830 17978 14854 17980
rect 14910 17978 14934 17980
rect 14772 17926 14774 17978
rect 14836 17926 14848 17978
rect 14910 17926 14912 17978
rect 14750 17924 14774 17926
rect 14830 17924 14854 17926
rect 14910 17924 14934 17926
rect 14694 17904 14990 17924
rect 14694 16892 14990 16912
rect 14750 16890 14774 16892
rect 14830 16890 14854 16892
rect 14910 16890 14934 16892
rect 14772 16838 14774 16890
rect 14836 16838 14848 16890
rect 14910 16838 14912 16890
rect 14750 16836 14774 16838
rect 14830 16836 14854 16838
rect 14910 16836 14934 16838
rect 14694 16816 14990 16836
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 14694 15804 14990 15824
rect 14750 15802 14774 15804
rect 14830 15802 14854 15804
rect 14910 15802 14934 15804
rect 14772 15750 14774 15802
rect 14836 15750 14848 15802
rect 14910 15750 14912 15802
rect 14750 15748 14774 15750
rect 14830 15748 14854 15750
rect 14910 15748 14934 15750
rect 14694 15728 14990 15748
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15856 15502 15884 15574
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15856 14958 15884 15438
rect 15948 14958 15976 15506
rect 16132 15366 16160 15982
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 14694 14716 14990 14736
rect 14750 14714 14774 14716
rect 14830 14714 14854 14716
rect 14910 14714 14934 14716
rect 14772 14662 14774 14714
rect 14836 14662 14848 14714
rect 14910 14662 14912 14714
rect 14750 14660 14774 14662
rect 14830 14660 14854 14662
rect 14910 14660 14934 14662
rect 14694 14640 14990 14660
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13360 13796 13412 13802
rect 13360 13738 13412 13744
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 11260 13084 11556 13104
rect 11316 13082 11340 13084
rect 11396 13082 11420 13084
rect 11476 13082 11500 13084
rect 11338 13030 11340 13082
rect 11402 13030 11414 13082
rect 11476 13030 11478 13082
rect 11316 13028 11340 13030
rect 11396 13028 11420 13030
rect 11476 13028 11500 13030
rect 11260 13008 11556 13028
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 11260 11996 11556 12016
rect 11316 11994 11340 11996
rect 11396 11994 11420 11996
rect 11476 11994 11500 11996
rect 11338 11942 11340 11994
rect 11402 11942 11414 11994
rect 11476 11942 11478 11994
rect 11316 11940 11340 11942
rect 11396 11940 11420 11942
rect 11476 11940 11500 11942
rect 11260 11920 11556 11940
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 7825 10364 8121 10384
rect 7881 10362 7905 10364
rect 7961 10362 7985 10364
rect 8041 10362 8065 10364
rect 7903 10310 7905 10362
rect 7967 10310 7979 10362
rect 8041 10310 8043 10362
rect 7881 10308 7905 10310
rect 7961 10308 7985 10310
rect 8041 10308 8065 10310
rect 7825 10288 8121 10308
rect 9968 9586 9996 10542
rect 10244 9602 10272 10542
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 10152 9574 10272 9602
rect 7825 9276 8121 9296
rect 7881 9274 7905 9276
rect 7961 9274 7985 9276
rect 8041 9274 8065 9276
rect 7903 9222 7905 9274
rect 7967 9222 7979 9274
rect 8041 9222 8043 9274
rect 7881 9220 7905 9222
rect 7961 9220 7985 9222
rect 8041 9220 8065 9222
rect 7825 9200 8121 9220
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7668 8090 7696 8978
rect 9968 8906 9996 9522
rect 10152 9518 10180 9574
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10428 9042 10456 11086
rect 10520 10810 10548 11630
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 7825 8188 8121 8208
rect 7881 8186 7905 8188
rect 7961 8186 7985 8188
rect 8041 8186 8065 8188
rect 7903 8134 7905 8186
rect 7967 8134 7979 8186
rect 8041 8134 8043 8186
rect 7881 8132 7905 8134
rect 7961 8132 7985 8134
rect 8041 8132 8065 8134
rect 7825 8112 8121 8132
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7300 6934 7328 7822
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7116 6186 7144 6802
rect 7300 6798 7328 6870
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7484 6322 7512 7686
rect 8680 7546 8708 8366
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7760 7206 7788 7346
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6012 4078 6040 4422
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 6104 3602 6132 4422
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 4390 3292 4686 3312
rect 4446 3290 4470 3292
rect 4526 3290 4550 3292
rect 4606 3290 4630 3292
rect 4468 3238 4470 3290
rect 4532 3238 4544 3290
rect 4606 3238 4608 3290
rect 4446 3236 4470 3238
rect 4526 3236 4550 3238
rect 4606 3236 4630 3238
rect 4390 3216 4686 3236
rect 4390 2204 4686 2224
rect 4446 2202 4470 2204
rect 4526 2202 4550 2204
rect 4606 2202 4630 2204
rect 4468 2150 4470 2202
rect 4532 2150 4544 2202
rect 4606 2150 4608 2202
rect 4446 2148 4470 2150
rect 4526 2148 4550 2150
rect 4606 2148 4630 2150
rect 4390 2128 4686 2148
rect 7116 800 7144 6122
rect 7668 5778 7696 6598
rect 7760 5914 7788 7142
rect 7825 7100 8121 7120
rect 7881 7098 7905 7100
rect 7961 7098 7985 7100
rect 8041 7098 8065 7100
rect 7903 7046 7905 7098
rect 7967 7046 7979 7098
rect 8041 7046 8043 7098
rect 7881 7044 7905 7046
rect 7961 7044 7985 7046
rect 8041 7044 8065 7046
rect 7825 7024 8121 7044
rect 8220 7002 8248 7278
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 7852 6322 7880 6870
rect 8772 6390 8800 8366
rect 9600 7342 9628 8774
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8864 7002 8892 7142
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 7825 6012 8121 6032
rect 7881 6010 7905 6012
rect 7961 6010 7985 6012
rect 8041 6010 8065 6012
rect 7903 5958 7905 6010
rect 7967 5958 7979 6010
rect 8041 5958 8043 6010
rect 7881 5956 7905 5958
rect 7961 5956 7985 5958
rect 8041 5956 8065 5958
rect 7825 5936 8121 5956
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7825 4924 8121 4944
rect 7881 4922 7905 4924
rect 7961 4922 7985 4924
rect 8041 4922 8065 4924
rect 7903 4870 7905 4922
rect 7967 4870 7979 4922
rect 8041 4870 8043 4922
rect 7881 4868 7905 4870
rect 7961 4868 7985 4870
rect 8041 4868 8065 4870
rect 7825 4848 8121 4868
rect 7825 3836 8121 3856
rect 7881 3834 7905 3836
rect 7961 3834 7985 3836
rect 8041 3834 8065 3836
rect 7903 3782 7905 3834
rect 7967 3782 7979 3834
rect 8041 3782 8043 3834
rect 7881 3780 7905 3782
rect 7961 3780 7985 3782
rect 8041 3780 8065 3782
rect 7825 3760 8121 3780
rect 7825 2748 8121 2768
rect 7881 2746 7905 2748
rect 7961 2746 7985 2748
rect 8041 2746 8065 2748
rect 7903 2694 7905 2746
rect 7967 2694 7979 2746
rect 8041 2694 8043 2746
rect 7881 2692 7905 2694
rect 7961 2692 7985 2694
rect 8041 2692 8065 2694
rect 7825 2672 8121 2692
rect 9968 800 9996 8842
rect 10428 6458 10456 8978
rect 10520 8974 10548 10474
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10612 8430 10640 11290
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11164 10266 11192 11154
rect 11260 10908 11556 10928
rect 11316 10906 11340 10908
rect 11396 10906 11420 10908
rect 11476 10906 11500 10908
rect 11338 10854 11340 10906
rect 11402 10854 11414 10906
rect 11476 10854 11478 10906
rect 11316 10852 11340 10854
rect 11396 10852 11420 10854
rect 11476 10852 11500 10854
rect 11260 10832 11556 10852
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11716 10130 11744 11494
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 10704 8634 10732 10066
rect 11164 9722 11192 10066
rect 11260 9820 11556 9840
rect 11316 9818 11340 9820
rect 11396 9818 11420 9820
rect 11476 9818 11500 9820
rect 11338 9766 11340 9818
rect 11402 9766 11414 9818
rect 11476 9766 11478 9818
rect 11316 9764 11340 9766
rect 11396 9764 11420 9766
rect 11476 9764 11500 9766
rect 11260 9744 11556 9764
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10796 9042 10824 9386
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 11260 8732 11556 8752
rect 11316 8730 11340 8732
rect 11396 8730 11420 8732
rect 11476 8730 11500 8732
rect 11338 8678 11340 8730
rect 11402 8678 11414 8730
rect 11476 8678 11478 8730
rect 11316 8676 11340 8678
rect 11396 8676 11420 8678
rect 11476 8676 11500 8678
rect 11260 8656 11556 8676
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 11260 7644 11556 7664
rect 11316 7642 11340 7644
rect 11396 7642 11420 7644
rect 11476 7642 11500 7644
rect 11338 7590 11340 7642
rect 11402 7590 11414 7642
rect 11476 7590 11478 7642
rect 11316 7588 11340 7590
rect 11396 7588 11420 7590
rect 11476 7588 11500 7590
rect 11260 7568 11556 7588
rect 11260 6556 11556 6576
rect 11316 6554 11340 6556
rect 11396 6554 11420 6556
rect 11476 6554 11500 6556
rect 11338 6502 11340 6554
rect 11402 6502 11414 6554
rect 11476 6502 11478 6554
rect 11316 6500 11340 6502
rect 11396 6500 11420 6502
rect 11476 6500 11500 6502
rect 11260 6480 11556 6500
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 11260 5468 11556 5488
rect 11316 5466 11340 5468
rect 11396 5466 11420 5468
rect 11476 5466 11500 5468
rect 11338 5414 11340 5466
rect 11402 5414 11414 5466
rect 11476 5414 11478 5466
rect 11316 5412 11340 5414
rect 11396 5412 11420 5414
rect 11476 5412 11500 5414
rect 11260 5392 11556 5412
rect 11260 4380 11556 4400
rect 11316 4378 11340 4380
rect 11396 4378 11420 4380
rect 11476 4378 11500 4380
rect 11338 4326 11340 4378
rect 11402 4326 11414 4378
rect 11476 4326 11478 4378
rect 11316 4324 11340 4326
rect 11396 4324 11420 4326
rect 11476 4324 11500 4326
rect 11260 4304 11556 4324
rect 11260 3292 11556 3312
rect 11316 3290 11340 3292
rect 11396 3290 11420 3292
rect 11476 3290 11500 3292
rect 11338 3238 11340 3290
rect 11402 3238 11414 3290
rect 11476 3238 11478 3290
rect 11316 3236 11340 3238
rect 11396 3236 11420 3238
rect 11476 3236 11500 3238
rect 11260 3216 11556 3236
rect 11260 2204 11556 2224
rect 11316 2202 11340 2204
rect 11396 2202 11420 2204
rect 11476 2202 11500 2204
rect 11338 2150 11340 2202
rect 11402 2150 11414 2202
rect 11476 2150 11478 2202
rect 11316 2148 11340 2150
rect 11396 2148 11420 2150
rect 11476 2148 11500 2150
rect 11260 2128 11556 2148
rect 12728 898 12756 12174
rect 13280 11234 13308 13330
rect 13372 13326 13400 13738
rect 13464 13394 13492 13806
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13464 12306 13492 13330
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13556 11898 13584 12718
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13648 11354 13676 13806
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13740 13394 13768 13670
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13740 12374 13768 13330
rect 14384 12782 14412 14214
rect 14568 14074 14596 14418
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14694 13628 14990 13648
rect 14750 13626 14774 13628
rect 14830 13626 14854 13628
rect 14910 13626 14934 13628
rect 14772 13574 14774 13626
rect 14836 13574 14848 13626
rect 14910 13574 14912 13626
rect 14750 13572 14774 13574
rect 14830 13572 14854 13574
rect 14910 13572 14934 13574
rect 14694 13552 14990 13572
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13832 11694 13860 12582
rect 14016 12374 14044 12718
rect 14694 12540 14990 12560
rect 14750 12538 14774 12540
rect 14830 12538 14854 12540
rect 14910 12538 14934 12540
rect 14772 12486 14774 12538
rect 14836 12486 14848 12538
rect 14910 12486 14912 12538
rect 14750 12484 14774 12486
rect 14830 12484 14854 12486
rect 14910 12484 14934 12486
rect 14694 12464 14990 12484
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 14694 11452 14990 11472
rect 14750 11450 14774 11452
rect 14830 11450 14854 11452
rect 14910 11450 14934 11452
rect 14772 11398 14774 11450
rect 14836 11398 14848 11450
rect 14910 11398 14912 11450
rect 14750 11396 14774 11398
rect 14830 11396 14854 11398
rect 14910 11396 14934 11398
rect 14694 11376 14990 11396
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13280 11218 13400 11234
rect 13280 11212 13412 11218
rect 13280 11206 13360 11212
rect 13360 11154 13412 11160
rect 13372 9178 13400 11154
rect 14694 10364 14990 10384
rect 14750 10362 14774 10364
rect 14830 10362 14854 10364
rect 14910 10362 14934 10364
rect 14772 10310 14774 10362
rect 14836 10310 14848 10362
rect 14910 10310 14912 10362
rect 14750 10308 14774 10310
rect 14830 10308 14854 10310
rect 14910 10308 14934 10310
rect 14694 10288 14990 10308
rect 14694 9276 14990 9296
rect 14750 9274 14774 9276
rect 14830 9274 14854 9276
rect 14910 9274 14934 9276
rect 14772 9222 14774 9274
rect 14836 9222 14848 9274
rect 14910 9222 14912 9274
rect 14750 9220 14774 9222
rect 14830 9220 14854 9222
rect 14910 9220 14934 9222
rect 14694 9200 14990 9220
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 14694 8188 14990 8208
rect 14750 8186 14774 8188
rect 14830 8186 14854 8188
rect 14910 8186 14934 8188
rect 14772 8134 14774 8186
rect 14836 8134 14848 8186
rect 14910 8134 14912 8186
rect 14750 8132 14774 8134
rect 14830 8132 14854 8134
rect 14910 8132 14934 8134
rect 14694 8112 14990 8132
rect 14694 7100 14990 7120
rect 14750 7098 14774 7100
rect 14830 7098 14854 7100
rect 14910 7098 14934 7100
rect 14772 7046 14774 7098
rect 14836 7046 14848 7098
rect 14910 7046 14912 7098
rect 14750 7044 14774 7046
rect 14830 7044 14854 7046
rect 14910 7044 14934 7046
rect 14694 7024 14990 7044
rect 14694 6012 14990 6032
rect 14750 6010 14774 6012
rect 14830 6010 14854 6012
rect 14910 6010 14934 6012
rect 14772 5958 14774 6010
rect 14836 5958 14848 6010
rect 14910 5958 14912 6010
rect 14750 5956 14774 5958
rect 14830 5956 14854 5958
rect 14910 5956 14934 5958
rect 14694 5936 14990 5956
rect 14694 4924 14990 4944
rect 14750 4922 14774 4924
rect 14830 4922 14854 4924
rect 14910 4922 14934 4924
rect 14772 4870 14774 4922
rect 14836 4870 14848 4922
rect 14910 4870 14912 4922
rect 14750 4868 14774 4870
rect 14830 4868 14854 4870
rect 14910 4868 14934 4870
rect 14694 4848 14990 4868
rect 14694 3836 14990 3856
rect 14750 3834 14774 3836
rect 14830 3834 14854 3836
rect 14910 3834 14934 3836
rect 14772 3782 14774 3834
rect 14836 3782 14848 3834
rect 14910 3782 14912 3834
rect 14750 3780 14774 3782
rect 14830 3780 14854 3782
rect 14910 3780 14934 3782
rect 14694 3760 14990 3780
rect 14694 2748 14990 2768
rect 14750 2746 14774 2748
rect 14830 2746 14854 2748
rect 14910 2746 14934 2748
rect 14772 2694 14774 2746
rect 14836 2694 14848 2746
rect 14910 2694 14912 2746
rect 14750 2692 14774 2694
rect 14830 2692 14854 2694
rect 14910 2692 14934 2694
rect 14694 2672 14990 2692
rect 15856 898 15884 14894
rect 16132 13530 16160 15302
rect 16224 15162 16252 16050
rect 16408 15706 16436 16050
rect 16500 16046 16528 24126
rect 18129 21788 18425 21808
rect 18185 21786 18209 21788
rect 18265 21786 18289 21788
rect 18345 21786 18369 21788
rect 18207 21734 18209 21786
rect 18271 21734 18283 21786
rect 18345 21734 18347 21786
rect 18185 21732 18209 21734
rect 18265 21732 18289 21734
rect 18345 21732 18369 21734
rect 18129 21712 18425 21732
rect 18129 20700 18425 20720
rect 18185 20698 18209 20700
rect 18265 20698 18289 20700
rect 18345 20698 18369 20700
rect 18207 20646 18209 20698
rect 18271 20646 18283 20698
rect 18345 20646 18347 20698
rect 18185 20644 18209 20646
rect 18265 20644 18289 20646
rect 18345 20644 18369 20646
rect 18129 20624 18425 20644
rect 18524 19802 18552 24202
rect 19062 23624 19118 23633
rect 19062 23559 19118 23568
rect 19076 21146 19104 23559
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19260 21010 19288 21490
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 19248 21004 19300 21010
rect 19248 20946 19300 20952
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 19892 21004 19944 21010
rect 19892 20946 19944 20952
rect 18524 19774 19012 19802
rect 18129 19612 18425 19632
rect 18185 19610 18209 19612
rect 18265 19610 18289 19612
rect 18345 19610 18369 19612
rect 18207 19558 18209 19610
rect 18271 19558 18283 19610
rect 18345 19558 18347 19610
rect 18185 19556 18209 19558
rect 18265 19556 18289 19558
rect 18345 19556 18369 19558
rect 18129 19536 18425 19556
rect 18984 19310 19012 19774
rect 18880 19304 18932 19310
rect 18880 19246 18932 19252
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18892 18698 18920 19246
rect 18984 18902 19012 19246
rect 19260 18970 19288 20946
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19536 19718 19564 20878
rect 19628 20330 19656 20946
rect 19904 20398 19932 20946
rect 20180 20534 20208 21422
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 20913 20484 21286
rect 21376 21010 21404 24202
rect 21364 21004 21416 21010
rect 21364 20946 21416 20952
rect 20442 20904 20498 20913
rect 20442 20839 20498 20848
rect 20168 20528 20220 20534
rect 20168 20470 20220 20476
rect 19892 20392 19944 20398
rect 19892 20334 19944 20340
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 19616 20324 19668 20330
rect 19616 20266 19668 20272
rect 19628 19922 19656 20266
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19904 19854 19932 20334
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18129 18524 18425 18544
rect 18185 18522 18209 18524
rect 18265 18522 18289 18524
rect 18345 18522 18369 18524
rect 18207 18470 18209 18522
rect 18271 18470 18283 18522
rect 18345 18470 18347 18522
rect 18185 18468 18209 18470
rect 18265 18468 18289 18470
rect 18345 18468 18369 18470
rect 18129 18448 18425 18468
rect 18892 18222 18920 18634
rect 18984 18290 19012 18838
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18129 17436 18425 17456
rect 18185 17434 18209 17436
rect 18265 17434 18289 17436
rect 18345 17434 18369 17436
rect 18207 17382 18209 17434
rect 18271 17382 18283 17434
rect 18345 17382 18347 17434
rect 18185 17380 18209 17382
rect 18265 17380 18289 17382
rect 18345 17380 18369 17382
rect 18129 17360 18425 17380
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16500 15586 16528 15982
rect 16408 15570 16528 15586
rect 17788 15570 17816 16730
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17880 15706 17908 16594
rect 18129 16348 18425 16368
rect 18185 16346 18209 16348
rect 18265 16346 18289 16348
rect 18345 16346 18369 16348
rect 18207 16294 18209 16346
rect 18271 16294 18283 16346
rect 18345 16294 18347 16346
rect 18185 16292 18209 16294
rect 18265 16292 18289 16294
rect 18345 16292 18369 16294
rect 18129 16272 18425 16292
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 16396 15564 16528 15570
rect 16448 15558 16528 15564
rect 17776 15564 17828 15570
rect 16396 15506 16448 15512
rect 17776 15506 17828 15512
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 18510 15328 18566 15337
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16592 14482 16620 14554
rect 16960 14482 16988 15302
rect 17052 14618 17080 15302
rect 18129 15260 18425 15280
rect 18510 15263 18566 15272
rect 18185 15258 18209 15260
rect 18265 15258 18289 15260
rect 18345 15258 18369 15260
rect 18207 15206 18209 15258
rect 18271 15206 18283 15258
rect 18345 15206 18347 15258
rect 18185 15204 18209 15206
rect 18265 15204 18289 15206
rect 18345 15204 18369 15206
rect 18129 15184 18425 15204
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17052 14482 17080 14554
rect 18524 14550 18552 15263
rect 18512 14544 18564 14550
rect 18512 14486 18564 14492
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 18129 14172 18425 14192
rect 18185 14170 18209 14172
rect 18265 14170 18289 14172
rect 18345 14170 18369 14172
rect 18207 14118 18209 14170
rect 18271 14118 18283 14170
rect 18345 14118 18347 14170
rect 18185 14116 18209 14118
rect 18265 14116 18289 14118
rect 18345 14116 18369 14118
rect 18129 14096 18425 14116
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 18129 13084 18425 13104
rect 18185 13082 18209 13084
rect 18265 13082 18289 13084
rect 18345 13082 18369 13084
rect 18207 13030 18209 13082
rect 18271 13030 18283 13082
rect 18345 13030 18347 13082
rect 18185 13028 18209 13030
rect 18265 13028 18289 13030
rect 18345 13028 18369 13030
rect 18129 13008 18425 13028
rect 18129 11996 18425 12016
rect 18185 11994 18209 11996
rect 18265 11994 18289 11996
rect 18345 11994 18369 11996
rect 18207 11942 18209 11994
rect 18271 11942 18283 11994
rect 18345 11942 18347 11994
rect 18185 11940 18209 11942
rect 18265 11940 18289 11942
rect 18345 11940 18369 11942
rect 18129 11920 18425 11940
rect 18129 10908 18425 10928
rect 18185 10906 18209 10908
rect 18265 10906 18289 10908
rect 18345 10906 18369 10908
rect 18207 10854 18209 10906
rect 18271 10854 18283 10906
rect 18345 10854 18347 10906
rect 18185 10852 18209 10854
rect 18265 10852 18289 10854
rect 18345 10852 18369 10854
rect 18129 10832 18425 10852
rect 18129 9820 18425 9840
rect 18185 9818 18209 9820
rect 18265 9818 18289 9820
rect 18345 9818 18369 9820
rect 18207 9766 18209 9818
rect 18271 9766 18283 9818
rect 18345 9766 18347 9818
rect 18185 9764 18209 9766
rect 18265 9764 18289 9766
rect 18345 9764 18369 9766
rect 18129 9744 18425 9764
rect 18129 8732 18425 8752
rect 18185 8730 18209 8732
rect 18265 8730 18289 8732
rect 18345 8730 18369 8732
rect 18207 8678 18209 8730
rect 18271 8678 18283 8730
rect 18345 8678 18347 8730
rect 18185 8676 18209 8678
rect 18265 8676 18289 8678
rect 18345 8676 18369 8678
rect 18129 8656 18425 8676
rect 18129 7644 18425 7664
rect 18185 7642 18209 7644
rect 18265 7642 18289 7644
rect 18345 7642 18369 7644
rect 18207 7590 18209 7642
rect 18271 7590 18283 7642
rect 18345 7590 18347 7642
rect 18185 7588 18209 7590
rect 18265 7588 18289 7590
rect 18345 7588 18369 7590
rect 18129 7568 18425 7588
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 18064 6905 18092 6938
rect 18050 6896 18106 6905
rect 18050 6831 18106 6840
rect 18129 6556 18425 6576
rect 18185 6554 18209 6556
rect 18265 6554 18289 6556
rect 18345 6554 18369 6556
rect 18207 6502 18209 6554
rect 18271 6502 18283 6554
rect 18345 6502 18347 6554
rect 18185 6500 18209 6502
rect 18265 6500 18289 6502
rect 18345 6500 18369 6502
rect 18129 6480 18425 6500
rect 18788 5636 18840 5642
rect 18788 5578 18840 5584
rect 18129 5468 18425 5488
rect 18185 5466 18209 5468
rect 18265 5466 18289 5468
rect 18345 5466 18369 5468
rect 18207 5414 18209 5466
rect 18271 5414 18283 5466
rect 18345 5414 18347 5466
rect 18185 5412 18209 5414
rect 18265 5412 18289 5414
rect 18345 5412 18369 5414
rect 18129 5392 18425 5412
rect 18129 4380 18425 4400
rect 18185 4378 18209 4380
rect 18265 4378 18289 4380
rect 18345 4378 18369 4380
rect 18207 4326 18209 4378
rect 18271 4326 18283 4378
rect 18345 4326 18347 4378
rect 18185 4324 18209 4326
rect 18265 4324 18289 4326
rect 18345 4324 18369 4326
rect 18129 4304 18425 4324
rect 18800 4185 18828 5578
rect 18786 4176 18842 4185
rect 18786 4111 18842 4120
rect 18129 3292 18425 3312
rect 18185 3290 18209 3292
rect 18265 3290 18289 3292
rect 18345 3290 18369 3292
rect 18207 3238 18209 3290
rect 18271 3238 18283 3290
rect 18345 3238 18347 3290
rect 18185 3236 18209 3238
rect 18265 3236 18289 3238
rect 18345 3236 18369 3238
rect 18129 3216 18425 3236
rect 18129 2204 18425 2224
rect 18185 2202 18209 2204
rect 18265 2202 18289 2204
rect 18345 2202 18369 2204
rect 18207 2150 18209 2202
rect 18271 2150 18283 2202
rect 18345 2150 18347 2202
rect 18185 2148 18209 2150
rect 18265 2148 18289 2150
rect 18345 2148 18369 2150
rect 18129 2128 18425 2148
rect 18892 898 18920 18158
rect 19260 17134 19288 18770
rect 19352 18766 19380 19178
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19890 18048 19946 18057
rect 19812 17746 19840 18022
rect 19890 17983 19946 17992
rect 19904 17814 19932 17983
rect 19892 17808 19944 17814
rect 19892 17750 19944 17756
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19352 17338 19380 17682
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 19260 16250 19288 17070
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19156 12708 19208 12714
rect 19156 12650 19208 12656
rect 19168 12481 19196 12650
rect 19154 12472 19210 12481
rect 19154 12407 19210 12416
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19260 9761 19288 9998
rect 19246 9752 19302 9761
rect 19246 9687 19302 9696
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 19260 1465 19288 2586
rect 19246 1456 19302 1465
rect 19246 1391 19302 1400
rect 20732 950 20760 20334
rect 12728 870 12848 898
rect 12820 800 12848 870
rect 15672 870 15884 898
rect 18524 870 18920 898
rect 20720 944 20772 950
rect 20720 886 20772 892
rect 21364 944 21416 950
rect 21364 886 21416 892
rect 15672 800 15700 870
rect 18524 800 18552 870
rect 21376 800 21404 886
rect 1398 0 1454 800
rect 4250 0 4306 800
rect 7102 0 7158 800
rect 9954 0 10010 800
rect 12806 0 12862 800
rect 15658 0 15714 800
rect 18510 0 18566 800
rect 21362 0 21418 800
<< via2 >>
rect 4390 21786 4446 21788
rect 4470 21786 4526 21788
rect 4550 21786 4606 21788
rect 4630 21786 4686 21788
rect 4390 21734 4416 21786
rect 4416 21734 4446 21786
rect 4470 21734 4480 21786
rect 4480 21734 4526 21786
rect 4550 21734 4596 21786
rect 4596 21734 4606 21786
rect 4630 21734 4660 21786
rect 4660 21734 4686 21786
rect 4390 21732 4446 21734
rect 4470 21732 4526 21734
rect 4550 21732 4606 21734
rect 4630 21732 4686 21734
rect 4390 20698 4446 20700
rect 4470 20698 4526 20700
rect 4550 20698 4606 20700
rect 4630 20698 4686 20700
rect 4390 20646 4416 20698
rect 4416 20646 4446 20698
rect 4470 20646 4480 20698
rect 4480 20646 4526 20698
rect 4550 20646 4596 20698
rect 4596 20646 4606 20698
rect 4630 20646 4660 20698
rect 4660 20646 4686 20698
rect 4390 20644 4446 20646
rect 4470 20644 4526 20646
rect 4550 20644 4606 20646
rect 4630 20644 4686 20646
rect 4390 19610 4446 19612
rect 4470 19610 4526 19612
rect 4550 19610 4606 19612
rect 4630 19610 4686 19612
rect 4390 19558 4416 19610
rect 4416 19558 4446 19610
rect 4470 19558 4480 19610
rect 4480 19558 4526 19610
rect 4550 19558 4596 19610
rect 4596 19558 4606 19610
rect 4630 19558 4660 19610
rect 4660 19558 4686 19610
rect 4390 19556 4446 19558
rect 4470 19556 4526 19558
rect 4550 19556 4606 19558
rect 4630 19556 4686 19558
rect 4390 18522 4446 18524
rect 4470 18522 4526 18524
rect 4550 18522 4606 18524
rect 4630 18522 4686 18524
rect 4390 18470 4416 18522
rect 4416 18470 4446 18522
rect 4470 18470 4480 18522
rect 4480 18470 4526 18522
rect 4550 18470 4596 18522
rect 4596 18470 4606 18522
rect 4630 18470 4660 18522
rect 4660 18470 4686 18522
rect 4390 18468 4446 18470
rect 4470 18468 4526 18470
rect 4550 18468 4606 18470
rect 4630 18468 4686 18470
rect 4390 17434 4446 17436
rect 4470 17434 4526 17436
rect 4550 17434 4606 17436
rect 4630 17434 4686 17436
rect 4390 17382 4416 17434
rect 4416 17382 4446 17434
rect 4470 17382 4480 17434
rect 4480 17382 4526 17434
rect 4550 17382 4596 17434
rect 4596 17382 4606 17434
rect 4630 17382 4660 17434
rect 4660 17382 4686 17434
rect 4390 17380 4446 17382
rect 4470 17380 4526 17382
rect 4550 17380 4606 17382
rect 4630 17380 4686 17382
rect 4390 16346 4446 16348
rect 4470 16346 4526 16348
rect 4550 16346 4606 16348
rect 4630 16346 4686 16348
rect 4390 16294 4416 16346
rect 4416 16294 4446 16346
rect 4470 16294 4480 16346
rect 4480 16294 4526 16346
rect 4550 16294 4596 16346
rect 4596 16294 4606 16346
rect 4630 16294 4660 16346
rect 4660 16294 4686 16346
rect 4390 16292 4446 16294
rect 4470 16292 4526 16294
rect 4550 16292 4606 16294
rect 4630 16292 4686 16294
rect 4390 15258 4446 15260
rect 4470 15258 4526 15260
rect 4550 15258 4606 15260
rect 4630 15258 4686 15260
rect 4390 15206 4416 15258
rect 4416 15206 4446 15258
rect 4470 15206 4480 15258
rect 4480 15206 4526 15258
rect 4550 15206 4596 15258
rect 4596 15206 4606 15258
rect 4630 15206 4660 15258
rect 4660 15206 4686 15258
rect 4390 15204 4446 15206
rect 4470 15204 4526 15206
rect 4550 15204 4606 15206
rect 4630 15204 4686 15206
rect 4390 14170 4446 14172
rect 4470 14170 4526 14172
rect 4550 14170 4606 14172
rect 4630 14170 4686 14172
rect 4390 14118 4416 14170
rect 4416 14118 4446 14170
rect 4470 14118 4480 14170
rect 4480 14118 4526 14170
rect 4550 14118 4596 14170
rect 4596 14118 4606 14170
rect 4630 14118 4660 14170
rect 4660 14118 4686 14170
rect 4390 14116 4446 14118
rect 4470 14116 4526 14118
rect 4550 14116 4606 14118
rect 4630 14116 4686 14118
rect 4390 13082 4446 13084
rect 4470 13082 4526 13084
rect 4550 13082 4606 13084
rect 4630 13082 4686 13084
rect 4390 13030 4416 13082
rect 4416 13030 4446 13082
rect 4470 13030 4480 13082
rect 4480 13030 4526 13082
rect 4550 13030 4596 13082
rect 4596 13030 4606 13082
rect 4630 13030 4660 13082
rect 4660 13030 4686 13082
rect 4390 13028 4446 13030
rect 4470 13028 4526 13030
rect 4550 13028 4606 13030
rect 4630 13028 4686 13030
rect 2870 12552 2926 12608
rect 4390 11994 4446 11996
rect 4470 11994 4526 11996
rect 4550 11994 4606 11996
rect 4630 11994 4686 11996
rect 4390 11942 4416 11994
rect 4416 11942 4446 11994
rect 4470 11942 4480 11994
rect 4480 11942 4526 11994
rect 4550 11942 4596 11994
rect 4596 11942 4606 11994
rect 4630 11942 4660 11994
rect 4660 11942 4686 11994
rect 4390 11940 4446 11942
rect 4470 11940 4526 11942
rect 4550 11940 4606 11942
rect 4630 11940 4686 11942
rect 4390 10906 4446 10908
rect 4470 10906 4526 10908
rect 4550 10906 4606 10908
rect 4630 10906 4686 10908
rect 4390 10854 4416 10906
rect 4416 10854 4446 10906
rect 4470 10854 4480 10906
rect 4480 10854 4526 10906
rect 4550 10854 4596 10906
rect 4596 10854 4606 10906
rect 4630 10854 4660 10906
rect 4660 10854 4686 10906
rect 4390 10852 4446 10854
rect 4470 10852 4526 10854
rect 4550 10852 4606 10854
rect 4630 10852 4686 10854
rect 4390 9818 4446 9820
rect 4470 9818 4526 9820
rect 4550 9818 4606 9820
rect 4630 9818 4686 9820
rect 4390 9766 4416 9818
rect 4416 9766 4446 9818
rect 4470 9766 4480 9818
rect 4480 9766 4526 9818
rect 4550 9766 4596 9818
rect 4596 9766 4606 9818
rect 4630 9766 4660 9818
rect 4660 9766 4686 9818
rect 4390 9764 4446 9766
rect 4470 9764 4526 9766
rect 4550 9764 4606 9766
rect 4630 9764 4686 9766
rect 4390 8730 4446 8732
rect 4470 8730 4526 8732
rect 4550 8730 4606 8732
rect 4630 8730 4686 8732
rect 4390 8678 4416 8730
rect 4416 8678 4446 8730
rect 4470 8678 4480 8730
rect 4480 8678 4526 8730
rect 4550 8678 4596 8730
rect 4596 8678 4606 8730
rect 4630 8678 4660 8730
rect 4660 8678 4686 8730
rect 4390 8676 4446 8678
rect 4470 8676 4526 8678
rect 4550 8676 4606 8678
rect 4630 8676 4686 8678
rect 4390 7642 4446 7644
rect 4470 7642 4526 7644
rect 4550 7642 4606 7644
rect 4630 7642 4686 7644
rect 4390 7590 4416 7642
rect 4416 7590 4446 7642
rect 4470 7590 4480 7642
rect 4480 7590 4526 7642
rect 4550 7590 4596 7642
rect 4596 7590 4606 7642
rect 4630 7590 4660 7642
rect 4660 7590 4686 7642
rect 4390 7588 4446 7590
rect 4470 7588 4526 7590
rect 4550 7588 4606 7590
rect 4630 7588 4686 7590
rect 4390 6554 4446 6556
rect 4470 6554 4526 6556
rect 4550 6554 4606 6556
rect 4630 6554 4686 6556
rect 4390 6502 4416 6554
rect 4416 6502 4446 6554
rect 4470 6502 4480 6554
rect 4480 6502 4526 6554
rect 4550 6502 4596 6554
rect 4596 6502 4606 6554
rect 4630 6502 4660 6554
rect 4660 6502 4686 6554
rect 4390 6500 4446 6502
rect 4470 6500 4526 6502
rect 4550 6500 4606 6502
rect 4630 6500 4686 6502
rect 4390 5466 4446 5468
rect 4470 5466 4526 5468
rect 4550 5466 4606 5468
rect 4630 5466 4686 5468
rect 4390 5414 4416 5466
rect 4416 5414 4446 5466
rect 4470 5414 4480 5466
rect 4480 5414 4526 5466
rect 4550 5414 4596 5466
rect 4596 5414 4606 5466
rect 4630 5414 4660 5466
rect 4660 5414 4686 5466
rect 4390 5412 4446 5414
rect 4470 5412 4526 5414
rect 4550 5412 4606 5414
rect 4630 5412 4686 5414
rect 4390 4378 4446 4380
rect 4470 4378 4526 4380
rect 4550 4378 4606 4380
rect 4630 4378 4686 4380
rect 4390 4326 4416 4378
rect 4416 4326 4446 4378
rect 4470 4326 4480 4378
rect 4480 4326 4526 4378
rect 4550 4326 4596 4378
rect 4596 4326 4606 4378
rect 4630 4326 4660 4378
rect 4660 4326 4686 4378
rect 4390 4324 4446 4326
rect 4470 4324 4526 4326
rect 4550 4324 4606 4326
rect 4630 4324 4686 4326
rect 7825 22330 7881 22332
rect 7905 22330 7961 22332
rect 7985 22330 8041 22332
rect 8065 22330 8121 22332
rect 7825 22278 7851 22330
rect 7851 22278 7881 22330
rect 7905 22278 7915 22330
rect 7915 22278 7961 22330
rect 7985 22278 8031 22330
rect 8031 22278 8041 22330
rect 8065 22278 8095 22330
rect 8095 22278 8121 22330
rect 7825 22276 7881 22278
rect 7905 22276 7961 22278
rect 7985 22276 8041 22278
rect 8065 22276 8121 22278
rect 7825 21242 7881 21244
rect 7905 21242 7961 21244
rect 7985 21242 8041 21244
rect 8065 21242 8121 21244
rect 7825 21190 7851 21242
rect 7851 21190 7881 21242
rect 7905 21190 7915 21242
rect 7915 21190 7961 21242
rect 7985 21190 8031 21242
rect 8031 21190 8041 21242
rect 8065 21190 8095 21242
rect 8095 21190 8121 21242
rect 7825 21188 7881 21190
rect 7905 21188 7961 21190
rect 7985 21188 8041 21190
rect 8065 21188 8121 21190
rect 7825 20154 7881 20156
rect 7905 20154 7961 20156
rect 7985 20154 8041 20156
rect 8065 20154 8121 20156
rect 7825 20102 7851 20154
rect 7851 20102 7881 20154
rect 7905 20102 7915 20154
rect 7915 20102 7961 20154
rect 7985 20102 8031 20154
rect 8031 20102 8041 20154
rect 8065 20102 8095 20154
rect 8095 20102 8121 20154
rect 7825 20100 7881 20102
rect 7905 20100 7961 20102
rect 7985 20100 8041 20102
rect 8065 20100 8121 20102
rect 7825 19066 7881 19068
rect 7905 19066 7961 19068
rect 7985 19066 8041 19068
rect 8065 19066 8121 19068
rect 7825 19014 7851 19066
rect 7851 19014 7881 19066
rect 7905 19014 7915 19066
rect 7915 19014 7961 19066
rect 7985 19014 8031 19066
rect 8031 19014 8041 19066
rect 8065 19014 8095 19066
rect 8095 19014 8121 19066
rect 7825 19012 7881 19014
rect 7905 19012 7961 19014
rect 7985 19012 8041 19014
rect 8065 19012 8121 19014
rect 7825 17978 7881 17980
rect 7905 17978 7961 17980
rect 7985 17978 8041 17980
rect 8065 17978 8121 17980
rect 7825 17926 7851 17978
rect 7851 17926 7881 17978
rect 7905 17926 7915 17978
rect 7915 17926 7961 17978
rect 7985 17926 8031 17978
rect 8031 17926 8041 17978
rect 8065 17926 8095 17978
rect 8095 17926 8121 17978
rect 7825 17924 7881 17926
rect 7905 17924 7961 17926
rect 7985 17924 8041 17926
rect 8065 17924 8121 17926
rect 7825 16890 7881 16892
rect 7905 16890 7961 16892
rect 7985 16890 8041 16892
rect 8065 16890 8121 16892
rect 7825 16838 7851 16890
rect 7851 16838 7881 16890
rect 7905 16838 7915 16890
rect 7915 16838 7961 16890
rect 7985 16838 8031 16890
rect 8031 16838 8041 16890
rect 8065 16838 8095 16890
rect 8095 16838 8121 16890
rect 7825 16836 7881 16838
rect 7905 16836 7961 16838
rect 7985 16836 8041 16838
rect 8065 16836 8121 16838
rect 7825 15802 7881 15804
rect 7905 15802 7961 15804
rect 7985 15802 8041 15804
rect 8065 15802 8121 15804
rect 7825 15750 7851 15802
rect 7851 15750 7881 15802
rect 7905 15750 7915 15802
rect 7915 15750 7961 15802
rect 7985 15750 8031 15802
rect 8031 15750 8041 15802
rect 8065 15750 8095 15802
rect 8095 15750 8121 15802
rect 7825 15748 7881 15750
rect 7905 15748 7961 15750
rect 7985 15748 8041 15750
rect 8065 15748 8121 15750
rect 7825 14714 7881 14716
rect 7905 14714 7961 14716
rect 7985 14714 8041 14716
rect 8065 14714 8121 14716
rect 7825 14662 7851 14714
rect 7851 14662 7881 14714
rect 7905 14662 7915 14714
rect 7915 14662 7961 14714
rect 7985 14662 8031 14714
rect 8031 14662 8041 14714
rect 8065 14662 8095 14714
rect 8095 14662 8121 14714
rect 7825 14660 7881 14662
rect 7905 14660 7961 14662
rect 7985 14660 8041 14662
rect 8065 14660 8121 14662
rect 7825 13626 7881 13628
rect 7905 13626 7961 13628
rect 7985 13626 8041 13628
rect 8065 13626 8121 13628
rect 7825 13574 7851 13626
rect 7851 13574 7881 13626
rect 7905 13574 7915 13626
rect 7915 13574 7961 13626
rect 7985 13574 8031 13626
rect 8031 13574 8041 13626
rect 8065 13574 8095 13626
rect 8095 13574 8121 13626
rect 7825 13572 7881 13574
rect 7905 13572 7961 13574
rect 7985 13572 8041 13574
rect 8065 13572 8121 13574
rect 7825 12538 7881 12540
rect 7905 12538 7961 12540
rect 7985 12538 8041 12540
rect 8065 12538 8121 12540
rect 7825 12486 7851 12538
rect 7851 12486 7881 12538
rect 7905 12486 7915 12538
rect 7915 12486 7961 12538
rect 7985 12486 8031 12538
rect 8031 12486 8041 12538
rect 8065 12486 8095 12538
rect 8095 12486 8121 12538
rect 7825 12484 7881 12486
rect 7905 12484 7961 12486
rect 7985 12484 8041 12486
rect 8065 12484 8121 12486
rect 7825 11450 7881 11452
rect 7905 11450 7961 11452
rect 7985 11450 8041 11452
rect 8065 11450 8121 11452
rect 7825 11398 7851 11450
rect 7851 11398 7881 11450
rect 7905 11398 7915 11450
rect 7915 11398 7961 11450
rect 7985 11398 8031 11450
rect 8031 11398 8041 11450
rect 8065 11398 8095 11450
rect 8095 11398 8121 11450
rect 7825 11396 7881 11398
rect 7905 11396 7961 11398
rect 7985 11396 8041 11398
rect 8065 11396 8121 11398
rect 11260 21786 11316 21788
rect 11340 21786 11396 21788
rect 11420 21786 11476 21788
rect 11500 21786 11556 21788
rect 11260 21734 11286 21786
rect 11286 21734 11316 21786
rect 11340 21734 11350 21786
rect 11350 21734 11396 21786
rect 11420 21734 11466 21786
rect 11466 21734 11476 21786
rect 11500 21734 11530 21786
rect 11530 21734 11556 21786
rect 11260 21732 11316 21734
rect 11340 21732 11396 21734
rect 11420 21732 11476 21734
rect 11500 21732 11556 21734
rect 11260 20698 11316 20700
rect 11340 20698 11396 20700
rect 11420 20698 11476 20700
rect 11500 20698 11556 20700
rect 11260 20646 11286 20698
rect 11286 20646 11316 20698
rect 11340 20646 11350 20698
rect 11350 20646 11396 20698
rect 11420 20646 11466 20698
rect 11466 20646 11476 20698
rect 11500 20646 11530 20698
rect 11530 20646 11556 20698
rect 11260 20644 11316 20646
rect 11340 20644 11396 20646
rect 11420 20644 11476 20646
rect 11500 20644 11556 20646
rect 11260 19610 11316 19612
rect 11340 19610 11396 19612
rect 11420 19610 11476 19612
rect 11500 19610 11556 19612
rect 11260 19558 11286 19610
rect 11286 19558 11316 19610
rect 11340 19558 11350 19610
rect 11350 19558 11396 19610
rect 11420 19558 11466 19610
rect 11466 19558 11476 19610
rect 11500 19558 11530 19610
rect 11530 19558 11556 19610
rect 11260 19556 11316 19558
rect 11340 19556 11396 19558
rect 11420 19556 11476 19558
rect 11500 19556 11556 19558
rect 11260 18522 11316 18524
rect 11340 18522 11396 18524
rect 11420 18522 11476 18524
rect 11500 18522 11556 18524
rect 11260 18470 11286 18522
rect 11286 18470 11316 18522
rect 11340 18470 11350 18522
rect 11350 18470 11396 18522
rect 11420 18470 11466 18522
rect 11466 18470 11476 18522
rect 11500 18470 11530 18522
rect 11530 18470 11556 18522
rect 11260 18468 11316 18470
rect 11340 18468 11396 18470
rect 11420 18468 11476 18470
rect 11500 18468 11556 18470
rect 11260 17434 11316 17436
rect 11340 17434 11396 17436
rect 11420 17434 11476 17436
rect 11500 17434 11556 17436
rect 11260 17382 11286 17434
rect 11286 17382 11316 17434
rect 11340 17382 11350 17434
rect 11350 17382 11396 17434
rect 11420 17382 11466 17434
rect 11466 17382 11476 17434
rect 11500 17382 11530 17434
rect 11530 17382 11556 17434
rect 11260 17380 11316 17382
rect 11340 17380 11396 17382
rect 11420 17380 11476 17382
rect 11500 17380 11556 17382
rect 11260 16346 11316 16348
rect 11340 16346 11396 16348
rect 11420 16346 11476 16348
rect 11500 16346 11556 16348
rect 11260 16294 11286 16346
rect 11286 16294 11316 16346
rect 11340 16294 11350 16346
rect 11350 16294 11396 16346
rect 11420 16294 11466 16346
rect 11466 16294 11476 16346
rect 11500 16294 11530 16346
rect 11530 16294 11556 16346
rect 11260 16292 11316 16294
rect 11340 16292 11396 16294
rect 11420 16292 11476 16294
rect 11500 16292 11556 16294
rect 11260 15258 11316 15260
rect 11340 15258 11396 15260
rect 11420 15258 11476 15260
rect 11500 15258 11556 15260
rect 11260 15206 11286 15258
rect 11286 15206 11316 15258
rect 11340 15206 11350 15258
rect 11350 15206 11396 15258
rect 11420 15206 11466 15258
rect 11466 15206 11476 15258
rect 11500 15206 11530 15258
rect 11530 15206 11556 15258
rect 11260 15204 11316 15206
rect 11340 15204 11396 15206
rect 11420 15204 11476 15206
rect 11500 15204 11556 15206
rect 11260 14170 11316 14172
rect 11340 14170 11396 14172
rect 11420 14170 11476 14172
rect 11500 14170 11556 14172
rect 11260 14118 11286 14170
rect 11286 14118 11316 14170
rect 11340 14118 11350 14170
rect 11350 14118 11396 14170
rect 11420 14118 11466 14170
rect 11466 14118 11476 14170
rect 11500 14118 11530 14170
rect 11530 14118 11556 14170
rect 11260 14116 11316 14118
rect 11340 14116 11396 14118
rect 11420 14116 11476 14118
rect 11500 14116 11556 14118
rect 14694 22330 14750 22332
rect 14774 22330 14830 22332
rect 14854 22330 14910 22332
rect 14934 22330 14990 22332
rect 14694 22278 14720 22330
rect 14720 22278 14750 22330
rect 14774 22278 14784 22330
rect 14784 22278 14830 22330
rect 14854 22278 14900 22330
rect 14900 22278 14910 22330
rect 14934 22278 14964 22330
rect 14964 22278 14990 22330
rect 14694 22276 14750 22278
rect 14774 22276 14830 22278
rect 14854 22276 14910 22278
rect 14934 22276 14990 22278
rect 14694 21242 14750 21244
rect 14774 21242 14830 21244
rect 14854 21242 14910 21244
rect 14934 21242 14990 21244
rect 14694 21190 14720 21242
rect 14720 21190 14750 21242
rect 14774 21190 14784 21242
rect 14784 21190 14830 21242
rect 14854 21190 14900 21242
rect 14900 21190 14910 21242
rect 14934 21190 14964 21242
rect 14964 21190 14990 21242
rect 14694 21188 14750 21190
rect 14774 21188 14830 21190
rect 14854 21188 14910 21190
rect 14934 21188 14990 21190
rect 14694 20154 14750 20156
rect 14774 20154 14830 20156
rect 14854 20154 14910 20156
rect 14934 20154 14990 20156
rect 14694 20102 14720 20154
rect 14720 20102 14750 20154
rect 14774 20102 14784 20154
rect 14784 20102 14830 20154
rect 14854 20102 14900 20154
rect 14900 20102 14910 20154
rect 14934 20102 14964 20154
rect 14964 20102 14990 20154
rect 14694 20100 14750 20102
rect 14774 20100 14830 20102
rect 14854 20100 14910 20102
rect 14934 20100 14990 20102
rect 14694 19066 14750 19068
rect 14774 19066 14830 19068
rect 14854 19066 14910 19068
rect 14934 19066 14990 19068
rect 14694 19014 14720 19066
rect 14720 19014 14750 19066
rect 14774 19014 14784 19066
rect 14784 19014 14830 19066
rect 14854 19014 14900 19066
rect 14900 19014 14910 19066
rect 14934 19014 14964 19066
rect 14964 19014 14990 19066
rect 14694 19012 14750 19014
rect 14774 19012 14830 19014
rect 14854 19012 14910 19014
rect 14934 19012 14990 19014
rect 14694 17978 14750 17980
rect 14774 17978 14830 17980
rect 14854 17978 14910 17980
rect 14934 17978 14990 17980
rect 14694 17926 14720 17978
rect 14720 17926 14750 17978
rect 14774 17926 14784 17978
rect 14784 17926 14830 17978
rect 14854 17926 14900 17978
rect 14900 17926 14910 17978
rect 14934 17926 14964 17978
rect 14964 17926 14990 17978
rect 14694 17924 14750 17926
rect 14774 17924 14830 17926
rect 14854 17924 14910 17926
rect 14934 17924 14990 17926
rect 14694 16890 14750 16892
rect 14774 16890 14830 16892
rect 14854 16890 14910 16892
rect 14934 16890 14990 16892
rect 14694 16838 14720 16890
rect 14720 16838 14750 16890
rect 14774 16838 14784 16890
rect 14784 16838 14830 16890
rect 14854 16838 14900 16890
rect 14900 16838 14910 16890
rect 14934 16838 14964 16890
rect 14964 16838 14990 16890
rect 14694 16836 14750 16838
rect 14774 16836 14830 16838
rect 14854 16836 14910 16838
rect 14934 16836 14990 16838
rect 14694 15802 14750 15804
rect 14774 15802 14830 15804
rect 14854 15802 14910 15804
rect 14934 15802 14990 15804
rect 14694 15750 14720 15802
rect 14720 15750 14750 15802
rect 14774 15750 14784 15802
rect 14784 15750 14830 15802
rect 14854 15750 14900 15802
rect 14900 15750 14910 15802
rect 14934 15750 14964 15802
rect 14964 15750 14990 15802
rect 14694 15748 14750 15750
rect 14774 15748 14830 15750
rect 14854 15748 14910 15750
rect 14934 15748 14990 15750
rect 14694 14714 14750 14716
rect 14774 14714 14830 14716
rect 14854 14714 14910 14716
rect 14934 14714 14990 14716
rect 14694 14662 14720 14714
rect 14720 14662 14750 14714
rect 14774 14662 14784 14714
rect 14784 14662 14830 14714
rect 14854 14662 14900 14714
rect 14900 14662 14910 14714
rect 14934 14662 14964 14714
rect 14964 14662 14990 14714
rect 14694 14660 14750 14662
rect 14774 14660 14830 14662
rect 14854 14660 14910 14662
rect 14934 14660 14990 14662
rect 11260 13082 11316 13084
rect 11340 13082 11396 13084
rect 11420 13082 11476 13084
rect 11500 13082 11556 13084
rect 11260 13030 11286 13082
rect 11286 13030 11316 13082
rect 11340 13030 11350 13082
rect 11350 13030 11396 13082
rect 11420 13030 11466 13082
rect 11466 13030 11476 13082
rect 11500 13030 11530 13082
rect 11530 13030 11556 13082
rect 11260 13028 11316 13030
rect 11340 13028 11396 13030
rect 11420 13028 11476 13030
rect 11500 13028 11556 13030
rect 11260 11994 11316 11996
rect 11340 11994 11396 11996
rect 11420 11994 11476 11996
rect 11500 11994 11556 11996
rect 11260 11942 11286 11994
rect 11286 11942 11316 11994
rect 11340 11942 11350 11994
rect 11350 11942 11396 11994
rect 11420 11942 11466 11994
rect 11466 11942 11476 11994
rect 11500 11942 11530 11994
rect 11530 11942 11556 11994
rect 11260 11940 11316 11942
rect 11340 11940 11396 11942
rect 11420 11940 11476 11942
rect 11500 11940 11556 11942
rect 7825 10362 7881 10364
rect 7905 10362 7961 10364
rect 7985 10362 8041 10364
rect 8065 10362 8121 10364
rect 7825 10310 7851 10362
rect 7851 10310 7881 10362
rect 7905 10310 7915 10362
rect 7915 10310 7961 10362
rect 7985 10310 8031 10362
rect 8031 10310 8041 10362
rect 8065 10310 8095 10362
rect 8095 10310 8121 10362
rect 7825 10308 7881 10310
rect 7905 10308 7961 10310
rect 7985 10308 8041 10310
rect 8065 10308 8121 10310
rect 7825 9274 7881 9276
rect 7905 9274 7961 9276
rect 7985 9274 8041 9276
rect 8065 9274 8121 9276
rect 7825 9222 7851 9274
rect 7851 9222 7881 9274
rect 7905 9222 7915 9274
rect 7915 9222 7961 9274
rect 7985 9222 8031 9274
rect 8031 9222 8041 9274
rect 8065 9222 8095 9274
rect 8095 9222 8121 9274
rect 7825 9220 7881 9222
rect 7905 9220 7961 9222
rect 7985 9220 8041 9222
rect 8065 9220 8121 9222
rect 7825 8186 7881 8188
rect 7905 8186 7961 8188
rect 7985 8186 8041 8188
rect 8065 8186 8121 8188
rect 7825 8134 7851 8186
rect 7851 8134 7881 8186
rect 7905 8134 7915 8186
rect 7915 8134 7961 8186
rect 7985 8134 8031 8186
rect 8031 8134 8041 8186
rect 8065 8134 8095 8186
rect 8095 8134 8121 8186
rect 7825 8132 7881 8134
rect 7905 8132 7961 8134
rect 7985 8132 8041 8134
rect 8065 8132 8121 8134
rect 4390 3290 4446 3292
rect 4470 3290 4526 3292
rect 4550 3290 4606 3292
rect 4630 3290 4686 3292
rect 4390 3238 4416 3290
rect 4416 3238 4446 3290
rect 4470 3238 4480 3290
rect 4480 3238 4526 3290
rect 4550 3238 4596 3290
rect 4596 3238 4606 3290
rect 4630 3238 4660 3290
rect 4660 3238 4686 3290
rect 4390 3236 4446 3238
rect 4470 3236 4526 3238
rect 4550 3236 4606 3238
rect 4630 3236 4686 3238
rect 4390 2202 4446 2204
rect 4470 2202 4526 2204
rect 4550 2202 4606 2204
rect 4630 2202 4686 2204
rect 4390 2150 4416 2202
rect 4416 2150 4446 2202
rect 4470 2150 4480 2202
rect 4480 2150 4526 2202
rect 4550 2150 4596 2202
rect 4596 2150 4606 2202
rect 4630 2150 4660 2202
rect 4660 2150 4686 2202
rect 4390 2148 4446 2150
rect 4470 2148 4526 2150
rect 4550 2148 4606 2150
rect 4630 2148 4686 2150
rect 7825 7098 7881 7100
rect 7905 7098 7961 7100
rect 7985 7098 8041 7100
rect 8065 7098 8121 7100
rect 7825 7046 7851 7098
rect 7851 7046 7881 7098
rect 7905 7046 7915 7098
rect 7915 7046 7961 7098
rect 7985 7046 8031 7098
rect 8031 7046 8041 7098
rect 8065 7046 8095 7098
rect 8095 7046 8121 7098
rect 7825 7044 7881 7046
rect 7905 7044 7961 7046
rect 7985 7044 8041 7046
rect 8065 7044 8121 7046
rect 7825 6010 7881 6012
rect 7905 6010 7961 6012
rect 7985 6010 8041 6012
rect 8065 6010 8121 6012
rect 7825 5958 7851 6010
rect 7851 5958 7881 6010
rect 7905 5958 7915 6010
rect 7915 5958 7961 6010
rect 7985 5958 8031 6010
rect 8031 5958 8041 6010
rect 8065 5958 8095 6010
rect 8095 5958 8121 6010
rect 7825 5956 7881 5958
rect 7905 5956 7961 5958
rect 7985 5956 8041 5958
rect 8065 5956 8121 5958
rect 7825 4922 7881 4924
rect 7905 4922 7961 4924
rect 7985 4922 8041 4924
rect 8065 4922 8121 4924
rect 7825 4870 7851 4922
rect 7851 4870 7881 4922
rect 7905 4870 7915 4922
rect 7915 4870 7961 4922
rect 7985 4870 8031 4922
rect 8031 4870 8041 4922
rect 8065 4870 8095 4922
rect 8095 4870 8121 4922
rect 7825 4868 7881 4870
rect 7905 4868 7961 4870
rect 7985 4868 8041 4870
rect 8065 4868 8121 4870
rect 7825 3834 7881 3836
rect 7905 3834 7961 3836
rect 7985 3834 8041 3836
rect 8065 3834 8121 3836
rect 7825 3782 7851 3834
rect 7851 3782 7881 3834
rect 7905 3782 7915 3834
rect 7915 3782 7961 3834
rect 7985 3782 8031 3834
rect 8031 3782 8041 3834
rect 8065 3782 8095 3834
rect 8095 3782 8121 3834
rect 7825 3780 7881 3782
rect 7905 3780 7961 3782
rect 7985 3780 8041 3782
rect 8065 3780 8121 3782
rect 7825 2746 7881 2748
rect 7905 2746 7961 2748
rect 7985 2746 8041 2748
rect 8065 2746 8121 2748
rect 7825 2694 7851 2746
rect 7851 2694 7881 2746
rect 7905 2694 7915 2746
rect 7915 2694 7961 2746
rect 7985 2694 8031 2746
rect 8031 2694 8041 2746
rect 8065 2694 8095 2746
rect 8095 2694 8121 2746
rect 7825 2692 7881 2694
rect 7905 2692 7961 2694
rect 7985 2692 8041 2694
rect 8065 2692 8121 2694
rect 11260 10906 11316 10908
rect 11340 10906 11396 10908
rect 11420 10906 11476 10908
rect 11500 10906 11556 10908
rect 11260 10854 11286 10906
rect 11286 10854 11316 10906
rect 11340 10854 11350 10906
rect 11350 10854 11396 10906
rect 11420 10854 11466 10906
rect 11466 10854 11476 10906
rect 11500 10854 11530 10906
rect 11530 10854 11556 10906
rect 11260 10852 11316 10854
rect 11340 10852 11396 10854
rect 11420 10852 11476 10854
rect 11500 10852 11556 10854
rect 11260 9818 11316 9820
rect 11340 9818 11396 9820
rect 11420 9818 11476 9820
rect 11500 9818 11556 9820
rect 11260 9766 11286 9818
rect 11286 9766 11316 9818
rect 11340 9766 11350 9818
rect 11350 9766 11396 9818
rect 11420 9766 11466 9818
rect 11466 9766 11476 9818
rect 11500 9766 11530 9818
rect 11530 9766 11556 9818
rect 11260 9764 11316 9766
rect 11340 9764 11396 9766
rect 11420 9764 11476 9766
rect 11500 9764 11556 9766
rect 11260 8730 11316 8732
rect 11340 8730 11396 8732
rect 11420 8730 11476 8732
rect 11500 8730 11556 8732
rect 11260 8678 11286 8730
rect 11286 8678 11316 8730
rect 11340 8678 11350 8730
rect 11350 8678 11396 8730
rect 11420 8678 11466 8730
rect 11466 8678 11476 8730
rect 11500 8678 11530 8730
rect 11530 8678 11556 8730
rect 11260 8676 11316 8678
rect 11340 8676 11396 8678
rect 11420 8676 11476 8678
rect 11500 8676 11556 8678
rect 11260 7642 11316 7644
rect 11340 7642 11396 7644
rect 11420 7642 11476 7644
rect 11500 7642 11556 7644
rect 11260 7590 11286 7642
rect 11286 7590 11316 7642
rect 11340 7590 11350 7642
rect 11350 7590 11396 7642
rect 11420 7590 11466 7642
rect 11466 7590 11476 7642
rect 11500 7590 11530 7642
rect 11530 7590 11556 7642
rect 11260 7588 11316 7590
rect 11340 7588 11396 7590
rect 11420 7588 11476 7590
rect 11500 7588 11556 7590
rect 11260 6554 11316 6556
rect 11340 6554 11396 6556
rect 11420 6554 11476 6556
rect 11500 6554 11556 6556
rect 11260 6502 11286 6554
rect 11286 6502 11316 6554
rect 11340 6502 11350 6554
rect 11350 6502 11396 6554
rect 11420 6502 11466 6554
rect 11466 6502 11476 6554
rect 11500 6502 11530 6554
rect 11530 6502 11556 6554
rect 11260 6500 11316 6502
rect 11340 6500 11396 6502
rect 11420 6500 11476 6502
rect 11500 6500 11556 6502
rect 11260 5466 11316 5468
rect 11340 5466 11396 5468
rect 11420 5466 11476 5468
rect 11500 5466 11556 5468
rect 11260 5414 11286 5466
rect 11286 5414 11316 5466
rect 11340 5414 11350 5466
rect 11350 5414 11396 5466
rect 11420 5414 11466 5466
rect 11466 5414 11476 5466
rect 11500 5414 11530 5466
rect 11530 5414 11556 5466
rect 11260 5412 11316 5414
rect 11340 5412 11396 5414
rect 11420 5412 11476 5414
rect 11500 5412 11556 5414
rect 11260 4378 11316 4380
rect 11340 4378 11396 4380
rect 11420 4378 11476 4380
rect 11500 4378 11556 4380
rect 11260 4326 11286 4378
rect 11286 4326 11316 4378
rect 11340 4326 11350 4378
rect 11350 4326 11396 4378
rect 11420 4326 11466 4378
rect 11466 4326 11476 4378
rect 11500 4326 11530 4378
rect 11530 4326 11556 4378
rect 11260 4324 11316 4326
rect 11340 4324 11396 4326
rect 11420 4324 11476 4326
rect 11500 4324 11556 4326
rect 11260 3290 11316 3292
rect 11340 3290 11396 3292
rect 11420 3290 11476 3292
rect 11500 3290 11556 3292
rect 11260 3238 11286 3290
rect 11286 3238 11316 3290
rect 11340 3238 11350 3290
rect 11350 3238 11396 3290
rect 11420 3238 11466 3290
rect 11466 3238 11476 3290
rect 11500 3238 11530 3290
rect 11530 3238 11556 3290
rect 11260 3236 11316 3238
rect 11340 3236 11396 3238
rect 11420 3236 11476 3238
rect 11500 3236 11556 3238
rect 11260 2202 11316 2204
rect 11340 2202 11396 2204
rect 11420 2202 11476 2204
rect 11500 2202 11556 2204
rect 11260 2150 11286 2202
rect 11286 2150 11316 2202
rect 11340 2150 11350 2202
rect 11350 2150 11396 2202
rect 11420 2150 11466 2202
rect 11466 2150 11476 2202
rect 11500 2150 11530 2202
rect 11530 2150 11556 2202
rect 11260 2148 11316 2150
rect 11340 2148 11396 2150
rect 11420 2148 11476 2150
rect 11500 2148 11556 2150
rect 14694 13626 14750 13628
rect 14774 13626 14830 13628
rect 14854 13626 14910 13628
rect 14934 13626 14990 13628
rect 14694 13574 14720 13626
rect 14720 13574 14750 13626
rect 14774 13574 14784 13626
rect 14784 13574 14830 13626
rect 14854 13574 14900 13626
rect 14900 13574 14910 13626
rect 14934 13574 14964 13626
rect 14964 13574 14990 13626
rect 14694 13572 14750 13574
rect 14774 13572 14830 13574
rect 14854 13572 14910 13574
rect 14934 13572 14990 13574
rect 14694 12538 14750 12540
rect 14774 12538 14830 12540
rect 14854 12538 14910 12540
rect 14934 12538 14990 12540
rect 14694 12486 14720 12538
rect 14720 12486 14750 12538
rect 14774 12486 14784 12538
rect 14784 12486 14830 12538
rect 14854 12486 14900 12538
rect 14900 12486 14910 12538
rect 14934 12486 14964 12538
rect 14964 12486 14990 12538
rect 14694 12484 14750 12486
rect 14774 12484 14830 12486
rect 14854 12484 14910 12486
rect 14934 12484 14990 12486
rect 14694 11450 14750 11452
rect 14774 11450 14830 11452
rect 14854 11450 14910 11452
rect 14934 11450 14990 11452
rect 14694 11398 14720 11450
rect 14720 11398 14750 11450
rect 14774 11398 14784 11450
rect 14784 11398 14830 11450
rect 14854 11398 14900 11450
rect 14900 11398 14910 11450
rect 14934 11398 14964 11450
rect 14964 11398 14990 11450
rect 14694 11396 14750 11398
rect 14774 11396 14830 11398
rect 14854 11396 14910 11398
rect 14934 11396 14990 11398
rect 14694 10362 14750 10364
rect 14774 10362 14830 10364
rect 14854 10362 14910 10364
rect 14934 10362 14990 10364
rect 14694 10310 14720 10362
rect 14720 10310 14750 10362
rect 14774 10310 14784 10362
rect 14784 10310 14830 10362
rect 14854 10310 14900 10362
rect 14900 10310 14910 10362
rect 14934 10310 14964 10362
rect 14964 10310 14990 10362
rect 14694 10308 14750 10310
rect 14774 10308 14830 10310
rect 14854 10308 14910 10310
rect 14934 10308 14990 10310
rect 14694 9274 14750 9276
rect 14774 9274 14830 9276
rect 14854 9274 14910 9276
rect 14934 9274 14990 9276
rect 14694 9222 14720 9274
rect 14720 9222 14750 9274
rect 14774 9222 14784 9274
rect 14784 9222 14830 9274
rect 14854 9222 14900 9274
rect 14900 9222 14910 9274
rect 14934 9222 14964 9274
rect 14964 9222 14990 9274
rect 14694 9220 14750 9222
rect 14774 9220 14830 9222
rect 14854 9220 14910 9222
rect 14934 9220 14990 9222
rect 14694 8186 14750 8188
rect 14774 8186 14830 8188
rect 14854 8186 14910 8188
rect 14934 8186 14990 8188
rect 14694 8134 14720 8186
rect 14720 8134 14750 8186
rect 14774 8134 14784 8186
rect 14784 8134 14830 8186
rect 14854 8134 14900 8186
rect 14900 8134 14910 8186
rect 14934 8134 14964 8186
rect 14964 8134 14990 8186
rect 14694 8132 14750 8134
rect 14774 8132 14830 8134
rect 14854 8132 14910 8134
rect 14934 8132 14990 8134
rect 14694 7098 14750 7100
rect 14774 7098 14830 7100
rect 14854 7098 14910 7100
rect 14934 7098 14990 7100
rect 14694 7046 14720 7098
rect 14720 7046 14750 7098
rect 14774 7046 14784 7098
rect 14784 7046 14830 7098
rect 14854 7046 14900 7098
rect 14900 7046 14910 7098
rect 14934 7046 14964 7098
rect 14964 7046 14990 7098
rect 14694 7044 14750 7046
rect 14774 7044 14830 7046
rect 14854 7044 14910 7046
rect 14934 7044 14990 7046
rect 14694 6010 14750 6012
rect 14774 6010 14830 6012
rect 14854 6010 14910 6012
rect 14934 6010 14990 6012
rect 14694 5958 14720 6010
rect 14720 5958 14750 6010
rect 14774 5958 14784 6010
rect 14784 5958 14830 6010
rect 14854 5958 14900 6010
rect 14900 5958 14910 6010
rect 14934 5958 14964 6010
rect 14964 5958 14990 6010
rect 14694 5956 14750 5958
rect 14774 5956 14830 5958
rect 14854 5956 14910 5958
rect 14934 5956 14990 5958
rect 14694 4922 14750 4924
rect 14774 4922 14830 4924
rect 14854 4922 14910 4924
rect 14934 4922 14990 4924
rect 14694 4870 14720 4922
rect 14720 4870 14750 4922
rect 14774 4870 14784 4922
rect 14784 4870 14830 4922
rect 14854 4870 14900 4922
rect 14900 4870 14910 4922
rect 14934 4870 14964 4922
rect 14964 4870 14990 4922
rect 14694 4868 14750 4870
rect 14774 4868 14830 4870
rect 14854 4868 14910 4870
rect 14934 4868 14990 4870
rect 14694 3834 14750 3836
rect 14774 3834 14830 3836
rect 14854 3834 14910 3836
rect 14934 3834 14990 3836
rect 14694 3782 14720 3834
rect 14720 3782 14750 3834
rect 14774 3782 14784 3834
rect 14784 3782 14830 3834
rect 14854 3782 14900 3834
rect 14900 3782 14910 3834
rect 14934 3782 14964 3834
rect 14964 3782 14990 3834
rect 14694 3780 14750 3782
rect 14774 3780 14830 3782
rect 14854 3780 14910 3782
rect 14934 3780 14990 3782
rect 14694 2746 14750 2748
rect 14774 2746 14830 2748
rect 14854 2746 14910 2748
rect 14934 2746 14990 2748
rect 14694 2694 14720 2746
rect 14720 2694 14750 2746
rect 14774 2694 14784 2746
rect 14784 2694 14830 2746
rect 14854 2694 14900 2746
rect 14900 2694 14910 2746
rect 14934 2694 14964 2746
rect 14964 2694 14990 2746
rect 14694 2692 14750 2694
rect 14774 2692 14830 2694
rect 14854 2692 14910 2694
rect 14934 2692 14990 2694
rect 18129 21786 18185 21788
rect 18209 21786 18265 21788
rect 18289 21786 18345 21788
rect 18369 21786 18425 21788
rect 18129 21734 18155 21786
rect 18155 21734 18185 21786
rect 18209 21734 18219 21786
rect 18219 21734 18265 21786
rect 18289 21734 18335 21786
rect 18335 21734 18345 21786
rect 18369 21734 18399 21786
rect 18399 21734 18425 21786
rect 18129 21732 18185 21734
rect 18209 21732 18265 21734
rect 18289 21732 18345 21734
rect 18369 21732 18425 21734
rect 18129 20698 18185 20700
rect 18209 20698 18265 20700
rect 18289 20698 18345 20700
rect 18369 20698 18425 20700
rect 18129 20646 18155 20698
rect 18155 20646 18185 20698
rect 18209 20646 18219 20698
rect 18219 20646 18265 20698
rect 18289 20646 18335 20698
rect 18335 20646 18345 20698
rect 18369 20646 18399 20698
rect 18399 20646 18425 20698
rect 18129 20644 18185 20646
rect 18209 20644 18265 20646
rect 18289 20644 18345 20646
rect 18369 20644 18425 20646
rect 19062 23568 19118 23624
rect 18129 19610 18185 19612
rect 18209 19610 18265 19612
rect 18289 19610 18345 19612
rect 18369 19610 18425 19612
rect 18129 19558 18155 19610
rect 18155 19558 18185 19610
rect 18209 19558 18219 19610
rect 18219 19558 18265 19610
rect 18289 19558 18335 19610
rect 18335 19558 18345 19610
rect 18369 19558 18399 19610
rect 18399 19558 18425 19610
rect 18129 19556 18185 19558
rect 18209 19556 18265 19558
rect 18289 19556 18345 19558
rect 18369 19556 18425 19558
rect 20442 20848 20498 20904
rect 18129 18522 18185 18524
rect 18209 18522 18265 18524
rect 18289 18522 18345 18524
rect 18369 18522 18425 18524
rect 18129 18470 18155 18522
rect 18155 18470 18185 18522
rect 18209 18470 18219 18522
rect 18219 18470 18265 18522
rect 18289 18470 18335 18522
rect 18335 18470 18345 18522
rect 18369 18470 18399 18522
rect 18399 18470 18425 18522
rect 18129 18468 18185 18470
rect 18209 18468 18265 18470
rect 18289 18468 18345 18470
rect 18369 18468 18425 18470
rect 18129 17434 18185 17436
rect 18209 17434 18265 17436
rect 18289 17434 18345 17436
rect 18369 17434 18425 17436
rect 18129 17382 18155 17434
rect 18155 17382 18185 17434
rect 18209 17382 18219 17434
rect 18219 17382 18265 17434
rect 18289 17382 18335 17434
rect 18335 17382 18345 17434
rect 18369 17382 18399 17434
rect 18399 17382 18425 17434
rect 18129 17380 18185 17382
rect 18209 17380 18265 17382
rect 18289 17380 18345 17382
rect 18369 17380 18425 17382
rect 18129 16346 18185 16348
rect 18209 16346 18265 16348
rect 18289 16346 18345 16348
rect 18369 16346 18425 16348
rect 18129 16294 18155 16346
rect 18155 16294 18185 16346
rect 18209 16294 18219 16346
rect 18219 16294 18265 16346
rect 18289 16294 18335 16346
rect 18335 16294 18345 16346
rect 18369 16294 18399 16346
rect 18399 16294 18425 16346
rect 18129 16292 18185 16294
rect 18209 16292 18265 16294
rect 18289 16292 18345 16294
rect 18369 16292 18425 16294
rect 18510 15272 18566 15328
rect 18129 15258 18185 15260
rect 18209 15258 18265 15260
rect 18289 15258 18345 15260
rect 18369 15258 18425 15260
rect 18129 15206 18155 15258
rect 18155 15206 18185 15258
rect 18209 15206 18219 15258
rect 18219 15206 18265 15258
rect 18289 15206 18335 15258
rect 18335 15206 18345 15258
rect 18369 15206 18399 15258
rect 18399 15206 18425 15258
rect 18129 15204 18185 15206
rect 18209 15204 18265 15206
rect 18289 15204 18345 15206
rect 18369 15204 18425 15206
rect 18129 14170 18185 14172
rect 18209 14170 18265 14172
rect 18289 14170 18345 14172
rect 18369 14170 18425 14172
rect 18129 14118 18155 14170
rect 18155 14118 18185 14170
rect 18209 14118 18219 14170
rect 18219 14118 18265 14170
rect 18289 14118 18335 14170
rect 18335 14118 18345 14170
rect 18369 14118 18399 14170
rect 18399 14118 18425 14170
rect 18129 14116 18185 14118
rect 18209 14116 18265 14118
rect 18289 14116 18345 14118
rect 18369 14116 18425 14118
rect 18129 13082 18185 13084
rect 18209 13082 18265 13084
rect 18289 13082 18345 13084
rect 18369 13082 18425 13084
rect 18129 13030 18155 13082
rect 18155 13030 18185 13082
rect 18209 13030 18219 13082
rect 18219 13030 18265 13082
rect 18289 13030 18335 13082
rect 18335 13030 18345 13082
rect 18369 13030 18399 13082
rect 18399 13030 18425 13082
rect 18129 13028 18185 13030
rect 18209 13028 18265 13030
rect 18289 13028 18345 13030
rect 18369 13028 18425 13030
rect 18129 11994 18185 11996
rect 18209 11994 18265 11996
rect 18289 11994 18345 11996
rect 18369 11994 18425 11996
rect 18129 11942 18155 11994
rect 18155 11942 18185 11994
rect 18209 11942 18219 11994
rect 18219 11942 18265 11994
rect 18289 11942 18335 11994
rect 18335 11942 18345 11994
rect 18369 11942 18399 11994
rect 18399 11942 18425 11994
rect 18129 11940 18185 11942
rect 18209 11940 18265 11942
rect 18289 11940 18345 11942
rect 18369 11940 18425 11942
rect 18129 10906 18185 10908
rect 18209 10906 18265 10908
rect 18289 10906 18345 10908
rect 18369 10906 18425 10908
rect 18129 10854 18155 10906
rect 18155 10854 18185 10906
rect 18209 10854 18219 10906
rect 18219 10854 18265 10906
rect 18289 10854 18335 10906
rect 18335 10854 18345 10906
rect 18369 10854 18399 10906
rect 18399 10854 18425 10906
rect 18129 10852 18185 10854
rect 18209 10852 18265 10854
rect 18289 10852 18345 10854
rect 18369 10852 18425 10854
rect 18129 9818 18185 9820
rect 18209 9818 18265 9820
rect 18289 9818 18345 9820
rect 18369 9818 18425 9820
rect 18129 9766 18155 9818
rect 18155 9766 18185 9818
rect 18209 9766 18219 9818
rect 18219 9766 18265 9818
rect 18289 9766 18335 9818
rect 18335 9766 18345 9818
rect 18369 9766 18399 9818
rect 18399 9766 18425 9818
rect 18129 9764 18185 9766
rect 18209 9764 18265 9766
rect 18289 9764 18345 9766
rect 18369 9764 18425 9766
rect 18129 8730 18185 8732
rect 18209 8730 18265 8732
rect 18289 8730 18345 8732
rect 18369 8730 18425 8732
rect 18129 8678 18155 8730
rect 18155 8678 18185 8730
rect 18209 8678 18219 8730
rect 18219 8678 18265 8730
rect 18289 8678 18335 8730
rect 18335 8678 18345 8730
rect 18369 8678 18399 8730
rect 18399 8678 18425 8730
rect 18129 8676 18185 8678
rect 18209 8676 18265 8678
rect 18289 8676 18345 8678
rect 18369 8676 18425 8678
rect 18129 7642 18185 7644
rect 18209 7642 18265 7644
rect 18289 7642 18345 7644
rect 18369 7642 18425 7644
rect 18129 7590 18155 7642
rect 18155 7590 18185 7642
rect 18209 7590 18219 7642
rect 18219 7590 18265 7642
rect 18289 7590 18335 7642
rect 18335 7590 18345 7642
rect 18369 7590 18399 7642
rect 18399 7590 18425 7642
rect 18129 7588 18185 7590
rect 18209 7588 18265 7590
rect 18289 7588 18345 7590
rect 18369 7588 18425 7590
rect 18050 6840 18106 6896
rect 18129 6554 18185 6556
rect 18209 6554 18265 6556
rect 18289 6554 18345 6556
rect 18369 6554 18425 6556
rect 18129 6502 18155 6554
rect 18155 6502 18185 6554
rect 18209 6502 18219 6554
rect 18219 6502 18265 6554
rect 18289 6502 18335 6554
rect 18335 6502 18345 6554
rect 18369 6502 18399 6554
rect 18399 6502 18425 6554
rect 18129 6500 18185 6502
rect 18209 6500 18265 6502
rect 18289 6500 18345 6502
rect 18369 6500 18425 6502
rect 18129 5466 18185 5468
rect 18209 5466 18265 5468
rect 18289 5466 18345 5468
rect 18369 5466 18425 5468
rect 18129 5414 18155 5466
rect 18155 5414 18185 5466
rect 18209 5414 18219 5466
rect 18219 5414 18265 5466
rect 18289 5414 18335 5466
rect 18335 5414 18345 5466
rect 18369 5414 18399 5466
rect 18399 5414 18425 5466
rect 18129 5412 18185 5414
rect 18209 5412 18265 5414
rect 18289 5412 18345 5414
rect 18369 5412 18425 5414
rect 18129 4378 18185 4380
rect 18209 4378 18265 4380
rect 18289 4378 18345 4380
rect 18369 4378 18425 4380
rect 18129 4326 18155 4378
rect 18155 4326 18185 4378
rect 18209 4326 18219 4378
rect 18219 4326 18265 4378
rect 18289 4326 18335 4378
rect 18335 4326 18345 4378
rect 18369 4326 18399 4378
rect 18399 4326 18425 4378
rect 18129 4324 18185 4326
rect 18209 4324 18265 4326
rect 18289 4324 18345 4326
rect 18369 4324 18425 4326
rect 18786 4120 18842 4176
rect 18129 3290 18185 3292
rect 18209 3290 18265 3292
rect 18289 3290 18345 3292
rect 18369 3290 18425 3292
rect 18129 3238 18155 3290
rect 18155 3238 18185 3290
rect 18209 3238 18219 3290
rect 18219 3238 18265 3290
rect 18289 3238 18335 3290
rect 18335 3238 18345 3290
rect 18369 3238 18399 3290
rect 18399 3238 18425 3290
rect 18129 3236 18185 3238
rect 18209 3236 18265 3238
rect 18289 3236 18345 3238
rect 18369 3236 18425 3238
rect 18129 2202 18185 2204
rect 18209 2202 18265 2204
rect 18289 2202 18345 2204
rect 18369 2202 18425 2204
rect 18129 2150 18155 2202
rect 18155 2150 18185 2202
rect 18209 2150 18219 2202
rect 18219 2150 18265 2202
rect 18289 2150 18335 2202
rect 18335 2150 18345 2202
rect 18369 2150 18399 2202
rect 18399 2150 18425 2202
rect 18129 2148 18185 2150
rect 18209 2148 18265 2150
rect 18289 2148 18345 2150
rect 18369 2148 18425 2150
rect 19890 17992 19946 18048
rect 19154 12416 19210 12472
rect 19246 9696 19302 9752
rect 19246 1400 19302 1456
<< metal3 >>
rect 19057 23626 19123 23629
rect 22058 23626 22858 23656
rect 19057 23624 22858 23626
rect 19057 23568 19062 23624
rect 19118 23568 22858 23624
rect 19057 23566 22858 23568
rect 19057 23563 19123 23566
rect 22058 23536 22858 23566
rect 7813 22336 8133 22337
rect 7813 22272 7821 22336
rect 7885 22272 7901 22336
rect 7965 22272 7981 22336
rect 8045 22272 8061 22336
rect 8125 22272 8133 22336
rect 7813 22271 8133 22272
rect 14682 22336 15002 22337
rect 14682 22272 14690 22336
rect 14754 22272 14770 22336
rect 14834 22272 14850 22336
rect 14914 22272 14930 22336
rect 14994 22272 15002 22336
rect 14682 22271 15002 22272
rect 4378 21792 4698 21793
rect 4378 21728 4386 21792
rect 4450 21728 4466 21792
rect 4530 21728 4546 21792
rect 4610 21728 4626 21792
rect 4690 21728 4698 21792
rect 4378 21727 4698 21728
rect 11248 21792 11568 21793
rect 11248 21728 11256 21792
rect 11320 21728 11336 21792
rect 11400 21728 11416 21792
rect 11480 21728 11496 21792
rect 11560 21728 11568 21792
rect 11248 21727 11568 21728
rect 18117 21792 18437 21793
rect 18117 21728 18125 21792
rect 18189 21728 18205 21792
rect 18269 21728 18285 21792
rect 18349 21728 18365 21792
rect 18429 21728 18437 21792
rect 18117 21727 18437 21728
rect 7813 21248 8133 21249
rect 7813 21184 7821 21248
rect 7885 21184 7901 21248
rect 7965 21184 7981 21248
rect 8045 21184 8061 21248
rect 8125 21184 8133 21248
rect 7813 21183 8133 21184
rect 14682 21248 15002 21249
rect 14682 21184 14690 21248
rect 14754 21184 14770 21248
rect 14834 21184 14850 21248
rect 14914 21184 14930 21248
rect 14994 21184 15002 21248
rect 14682 21183 15002 21184
rect 20437 20906 20503 20909
rect 22058 20906 22858 20936
rect 20437 20904 22858 20906
rect 20437 20848 20442 20904
rect 20498 20848 22858 20904
rect 20437 20846 22858 20848
rect 20437 20843 20503 20846
rect 22058 20816 22858 20846
rect 4378 20704 4698 20705
rect 4378 20640 4386 20704
rect 4450 20640 4466 20704
rect 4530 20640 4546 20704
rect 4610 20640 4626 20704
rect 4690 20640 4698 20704
rect 4378 20639 4698 20640
rect 11248 20704 11568 20705
rect 11248 20640 11256 20704
rect 11320 20640 11336 20704
rect 11400 20640 11416 20704
rect 11480 20640 11496 20704
rect 11560 20640 11568 20704
rect 11248 20639 11568 20640
rect 18117 20704 18437 20705
rect 18117 20640 18125 20704
rect 18189 20640 18205 20704
rect 18269 20640 18285 20704
rect 18349 20640 18365 20704
rect 18429 20640 18437 20704
rect 18117 20639 18437 20640
rect 7813 20160 8133 20161
rect 7813 20096 7821 20160
rect 7885 20096 7901 20160
rect 7965 20096 7981 20160
rect 8045 20096 8061 20160
rect 8125 20096 8133 20160
rect 7813 20095 8133 20096
rect 14682 20160 15002 20161
rect 14682 20096 14690 20160
rect 14754 20096 14770 20160
rect 14834 20096 14850 20160
rect 14914 20096 14930 20160
rect 14994 20096 15002 20160
rect 14682 20095 15002 20096
rect 4378 19616 4698 19617
rect 4378 19552 4386 19616
rect 4450 19552 4466 19616
rect 4530 19552 4546 19616
rect 4610 19552 4626 19616
rect 4690 19552 4698 19616
rect 4378 19551 4698 19552
rect 11248 19616 11568 19617
rect 11248 19552 11256 19616
rect 11320 19552 11336 19616
rect 11400 19552 11416 19616
rect 11480 19552 11496 19616
rect 11560 19552 11568 19616
rect 11248 19551 11568 19552
rect 18117 19616 18437 19617
rect 18117 19552 18125 19616
rect 18189 19552 18205 19616
rect 18269 19552 18285 19616
rect 18349 19552 18365 19616
rect 18429 19552 18437 19616
rect 18117 19551 18437 19552
rect 7813 19072 8133 19073
rect 7813 19008 7821 19072
rect 7885 19008 7901 19072
rect 7965 19008 7981 19072
rect 8045 19008 8061 19072
rect 8125 19008 8133 19072
rect 7813 19007 8133 19008
rect 14682 19072 15002 19073
rect 14682 19008 14690 19072
rect 14754 19008 14770 19072
rect 14834 19008 14850 19072
rect 14914 19008 14930 19072
rect 14994 19008 15002 19072
rect 14682 19007 15002 19008
rect 4378 18528 4698 18529
rect 4378 18464 4386 18528
rect 4450 18464 4466 18528
rect 4530 18464 4546 18528
rect 4610 18464 4626 18528
rect 4690 18464 4698 18528
rect 4378 18463 4698 18464
rect 11248 18528 11568 18529
rect 11248 18464 11256 18528
rect 11320 18464 11336 18528
rect 11400 18464 11416 18528
rect 11480 18464 11496 18528
rect 11560 18464 11568 18528
rect 11248 18463 11568 18464
rect 18117 18528 18437 18529
rect 18117 18464 18125 18528
rect 18189 18464 18205 18528
rect 18269 18464 18285 18528
rect 18349 18464 18365 18528
rect 18429 18464 18437 18528
rect 18117 18463 18437 18464
rect 19885 18050 19951 18053
rect 22058 18050 22858 18080
rect 19885 18048 22858 18050
rect 19885 17992 19890 18048
rect 19946 17992 22858 18048
rect 19885 17990 22858 17992
rect 19885 17987 19951 17990
rect 7813 17984 8133 17985
rect 7813 17920 7821 17984
rect 7885 17920 7901 17984
rect 7965 17920 7981 17984
rect 8045 17920 8061 17984
rect 8125 17920 8133 17984
rect 7813 17919 8133 17920
rect 14682 17984 15002 17985
rect 14682 17920 14690 17984
rect 14754 17920 14770 17984
rect 14834 17920 14850 17984
rect 14914 17920 14930 17984
rect 14994 17920 15002 17984
rect 22058 17960 22858 17990
rect 14682 17919 15002 17920
rect 4378 17440 4698 17441
rect 4378 17376 4386 17440
rect 4450 17376 4466 17440
rect 4530 17376 4546 17440
rect 4610 17376 4626 17440
rect 4690 17376 4698 17440
rect 4378 17375 4698 17376
rect 11248 17440 11568 17441
rect 11248 17376 11256 17440
rect 11320 17376 11336 17440
rect 11400 17376 11416 17440
rect 11480 17376 11496 17440
rect 11560 17376 11568 17440
rect 11248 17375 11568 17376
rect 18117 17440 18437 17441
rect 18117 17376 18125 17440
rect 18189 17376 18205 17440
rect 18269 17376 18285 17440
rect 18349 17376 18365 17440
rect 18429 17376 18437 17440
rect 18117 17375 18437 17376
rect 7813 16896 8133 16897
rect 7813 16832 7821 16896
rect 7885 16832 7901 16896
rect 7965 16832 7981 16896
rect 8045 16832 8061 16896
rect 8125 16832 8133 16896
rect 7813 16831 8133 16832
rect 14682 16896 15002 16897
rect 14682 16832 14690 16896
rect 14754 16832 14770 16896
rect 14834 16832 14850 16896
rect 14914 16832 14930 16896
rect 14994 16832 15002 16896
rect 14682 16831 15002 16832
rect 4378 16352 4698 16353
rect 4378 16288 4386 16352
rect 4450 16288 4466 16352
rect 4530 16288 4546 16352
rect 4610 16288 4626 16352
rect 4690 16288 4698 16352
rect 4378 16287 4698 16288
rect 11248 16352 11568 16353
rect 11248 16288 11256 16352
rect 11320 16288 11336 16352
rect 11400 16288 11416 16352
rect 11480 16288 11496 16352
rect 11560 16288 11568 16352
rect 11248 16287 11568 16288
rect 18117 16352 18437 16353
rect 18117 16288 18125 16352
rect 18189 16288 18205 16352
rect 18269 16288 18285 16352
rect 18349 16288 18365 16352
rect 18429 16288 18437 16352
rect 18117 16287 18437 16288
rect 7813 15808 8133 15809
rect 7813 15744 7821 15808
rect 7885 15744 7901 15808
rect 7965 15744 7981 15808
rect 8045 15744 8061 15808
rect 8125 15744 8133 15808
rect 7813 15743 8133 15744
rect 14682 15808 15002 15809
rect 14682 15744 14690 15808
rect 14754 15744 14770 15808
rect 14834 15744 14850 15808
rect 14914 15744 14930 15808
rect 14994 15744 15002 15808
rect 14682 15743 15002 15744
rect 18505 15330 18571 15333
rect 22058 15330 22858 15360
rect 18505 15328 22858 15330
rect 18505 15272 18510 15328
rect 18566 15272 22858 15328
rect 18505 15270 22858 15272
rect 18505 15267 18571 15270
rect 4378 15264 4698 15265
rect 4378 15200 4386 15264
rect 4450 15200 4466 15264
rect 4530 15200 4546 15264
rect 4610 15200 4626 15264
rect 4690 15200 4698 15264
rect 4378 15199 4698 15200
rect 11248 15264 11568 15265
rect 11248 15200 11256 15264
rect 11320 15200 11336 15264
rect 11400 15200 11416 15264
rect 11480 15200 11496 15264
rect 11560 15200 11568 15264
rect 11248 15199 11568 15200
rect 18117 15264 18437 15265
rect 18117 15200 18125 15264
rect 18189 15200 18205 15264
rect 18269 15200 18285 15264
rect 18349 15200 18365 15264
rect 18429 15200 18437 15264
rect 22058 15240 22858 15270
rect 18117 15199 18437 15200
rect 7813 14720 8133 14721
rect 7813 14656 7821 14720
rect 7885 14656 7901 14720
rect 7965 14656 7981 14720
rect 8045 14656 8061 14720
rect 8125 14656 8133 14720
rect 7813 14655 8133 14656
rect 14682 14720 15002 14721
rect 14682 14656 14690 14720
rect 14754 14656 14770 14720
rect 14834 14656 14850 14720
rect 14914 14656 14930 14720
rect 14994 14656 15002 14720
rect 14682 14655 15002 14656
rect 4378 14176 4698 14177
rect 4378 14112 4386 14176
rect 4450 14112 4466 14176
rect 4530 14112 4546 14176
rect 4610 14112 4626 14176
rect 4690 14112 4698 14176
rect 4378 14111 4698 14112
rect 11248 14176 11568 14177
rect 11248 14112 11256 14176
rect 11320 14112 11336 14176
rect 11400 14112 11416 14176
rect 11480 14112 11496 14176
rect 11560 14112 11568 14176
rect 11248 14111 11568 14112
rect 18117 14176 18437 14177
rect 18117 14112 18125 14176
rect 18189 14112 18205 14176
rect 18269 14112 18285 14176
rect 18349 14112 18365 14176
rect 18429 14112 18437 14176
rect 18117 14111 18437 14112
rect 7813 13632 8133 13633
rect 7813 13568 7821 13632
rect 7885 13568 7901 13632
rect 7965 13568 7981 13632
rect 8045 13568 8061 13632
rect 8125 13568 8133 13632
rect 7813 13567 8133 13568
rect 14682 13632 15002 13633
rect 14682 13568 14690 13632
rect 14754 13568 14770 13632
rect 14834 13568 14850 13632
rect 14914 13568 14930 13632
rect 14994 13568 15002 13632
rect 14682 13567 15002 13568
rect 4378 13088 4698 13089
rect 4378 13024 4386 13088
rect 4450 13024 4466 13088
rect 4530 13024 4546 13088
rect 4610 13024 4626 13088
rect 4690 13024 4698 13088
rect 4378 13023 4698 13024
rect 11248 13088 11568 13089
rect 11248 13024 11256 13088
rect 11320 13024 11336 13088
rect 11400 13024 11416 13088
rect 11480 13024 11496 13088
rect 11560 13024 11568 13088
rect 11248 13023 11568 13024
rect 18117 13088 18437 13089
rect 18117 13024 18125 13088
rect 18189 13024 18205 13088
rect 18269 13024 18285 13088
rect 18349 13024 18365 13088
rect 18429 13024 18437 13088
rect 18117 13023 18437 13024
rect 0 12610 800 12640
rect 2865 12610 2931 12613
rect 0 12608 2931 12610
rect 0 12552 2870 12608
rect 2926 12552 2931 12608
rect 0 12550 2931 12552
rect 0 12520 800 12550
rect 2865 12547 2931 12550
rect 7813 12544 8133 12545
rect 7813 12480 7821 12544
rect 7885 12480 7901 12544
rect 7965 12480 7981 12544
rect 8045 12480 8061 12544
rect 8125 12480 8133 12544
rect 7813 12479 8133 12480
rect 14682 12544 15002 12545
rect 14682 12480 14690 12544
rect 14754 12480 14770 12544
rect 14834 12480 14850 12544
rect 14914 12480 14930 12544
rect 14994 12480 15002 12544
rect 14682 12479 15002 12480
rect 19149 12474 19215 12477
rect 22058 12474 22858 12504
rect 19149 12472 22858 12474
rect 19149 12416 19154 12472
rect 19210 12416 22858 12472
rect 19149 12414 22858 12416
rect 19149 12411 19215 12414
rect 22058 12384 22858 12414
rect 4378 12000 4698 12001
rect 4378 11936 4386 12000
rect 4450 11936 4466 12000
rect 4530 11936 4546 12000
rect 4610 11936 4626 12000
rect 4690 11936 4698 12000
rect 4378 11935 4698 11936
rect 11248 12000 11568 12001
rect 11248 11936 11256 12000
rect 11320 11936 11336 12000
rect 11400 11936 11416 12000
rect 11480 11936 11496 12000
rect 11560 11936 11568 12000
rect 11248 11935 11568 11936
rect 18117 12000 18437 12001
rect 18117 11936 18125 12000
rect 18189 11936 18205 12000
rect 18269 11936 18285 12000
rect 18349 11936 18365 12000
rect 18429 11936 18437 12000
rect 18117 11935 18437 11936
rect 7813 11456 8133 11457
rect 7813 11392 7821 11456
rect 7885 11392 7901 11456
rect 7965 11392 7981 11456
rect 8045 11392 8061 11456
rect 8125 11392 8133 11456
rect 7813 11391 8133 11392
rect 14682 11456 15002 11457
rect 14682 11392 14690 11456
rect 14754 11392 14770 11456
rect 14834 11392 14850 11456
rect 14914 11392 14930 11456
rect 14994 11392 15002 11456
rect 14682 11391 15002 11392
rect 4378 10912 4698 10913
rect 4378 10848 4386 10912
rect 4450 10848 4466 10912
rect 4530 10848 4546 10912
rect 4610 10848 4626 10912
rect 4690 10848 4698 10912
rect 4378 10847 4698 10848
rect 11248 10912 11568 10913
rect 11248 10848 11256 10912
rect 11320 10848 11336 10912
rect 11400 10848 11416 10912
rect 11480 10848 11496 10912
rect 11560 10848 11568 10912
rect 11248 10847 11568 10848
rect 18117 10912 18437 10913
rect 18117 10848 18125 10912
rect 18189 10848 18205 10912
rect 18269 10848 18285 10912
rect 18349 10848 18365 10912
rect 18429 10848 18437 10912
rect 18117 10847 18437 10848
rect 7813 10368 8133 10369
rect 7813 10304 7821 10368
rect 7885 10304 7901 10368
rect 7965 10304 7981 10368
rect 8045 10304 8061 10368
rect 8125 10304 8133 10368
rect 7813 10303 8133 10304
rect 14682 10368 15002 10369
rect 14682 10304 14690 10368
rect 14754 10304 14770 10368
rect 14834 10304 14850 10368
rect 14914 10304 14930 10368
rect 14994 10304 15002 10368
rect 14682 10303 15002 10304
rect 4378 9824 4698 9825
rect 4378 9760 4386 9824
rect 4450 9760 4466 9824
rect 4530 9760 4546 9824
rect 4610 9760 4626 9824
rect 4690 9760 4698 9824
rect 4378 9759 4698 9760
rect 11248 9824 11568 9825
rect 11248 9760 11256 9824
rect 11320 9760 11336 9824
rect 11400 9760 11416 9824
rect 11480 9760 11496 9824
rect 11560 9760 11568 9824
rect 11248 9759 11568 9760
rect 18117 9824 18437 9825
rect 18117 9760 18125 9824
rect 18189 9760 18205 9824
rect 18269 9760 18285 9824
rect 18349 9760 18365 9824
rect 18429 9760 18437 9824
rect 18117 9759 18437 9760
rect 19241 9754 19307 9757
rect 22058 9754 22858 9784
rect 19241 9752 22858 9754
rect 19241 9696 19246 9752
rect 19302 9696 22858 9752
rect 19241 9694 22858 9696
rect 19241 9691 19307 9694
rect 22058 9664 22858 9694
rect 7813 9280 8133 9281
rect 7813 9216 7821 9280
rect 7885 9216 7901 9280
rect 7965 9216 7981 9280
rect 8045 9216 8061 9280
rect 8125 9216 8133 9280
rect 7813 9215 8133 9216
rect 14682 9280 15002 9281
rect 14682 9216 14690 9280
rect 14754 9216 14770 9280
rect 14834 9216 14850 9280
rect 14914 9216 14930 9280
rect 14994 9216 15002 9280
rect 14682 9215 15002 9216
rect 4378 8736 4698 8737
rect 4378 8672 4386 8736
rect 4450 8672 4466 8736
rect 4530 8672 4546 8736
rect 4610 8672 4626 8736
rect 4690 8672 4698 8736
rect 4378 8671 4698 8672
rect 11248 8736 11568 8737
rect 11248 8672 11256 8736
rect 11320 8672 11336 8736
rect 11400 8672 11416 8736
rect 11480 8672 11496 8736
rect 11560 8672 11568 8736
rect 11248 8671 11568 8672
rect 18117 8736 18437 8737
rect 18117 8672 18125 8736
rect 18189 8672 18205 8736
rect 18269 8672 18285 8736
rect 18349 8672 18365 8736
rect 18429 8672 18437 8736
rect 18117 8671 18437 8672
rect 7813 8192 8133 8193
rect 7813 8128 7821 8192
rect 7885 8128 7901 8192
rect 7965 8128 7981 8192
rect 8045 8128 8061 8192
rect 8125 8128 8133 8192
rect 7813 8127 8133 8128
rect 14682 8192 15002 8193
rect 14682 8128 14690 8192
rect 14754 8128 14770 8192
rect 14834 8128 14850 8192
rect 14914 8128 14930 8192
rect 14994 8128 15002 8192
rect 14682 8127 15002 8128
rect 4378 7648 4698 7649
rect 4378 7584 4386 7648
rect 4450 7584 4466 7648
rect 4530 7584 4546 7648
rect 4610 7584 4626 7648
rect 4690 7584 4698 7648
rect 4378 7583 4698 7584
rect 11248 7648 11568 7649
rect 11248 7584 11256 7648
rect 11320 7584 11336 7648
rect 11400 7584 11416 7648
rect 11480 7584 11496 7648
rect 11560 7584 11568 7648
rect 11248 7583 11568 7584
rect 18117 7648 18437 7649
rect 18117 7584 18125 7648
rect 18189 7584 18205 7648
rect 18269 7584 18285 7648
rect 18349 7584 18365 7648
rect 18429 7584 18437 7648
rect 18117 7583 18437 7584
rect 7813 7104 8133 7105
rect 7813 7040 7821 7104
rect 7885 7040 7901 7104
rect 7965 7040 7981 7104
rect 8045 7040 8061 7104
rect 8125 7040 8133 7104
rect 7813 7039 8133 7040
rect 14682 7104 15002 7105
rect 14682 7040 14690 7104
rect 14754 7040 14770 7104
rect 14834 7040 14850 7104
rect 14914 7040 14930 7104
rect 14994 7040 15002 7104
rect 14682 7039 15002 7040
rect 18045 6898 18111 6901
rect 22058 6898 22858 6928
rect 18045 6896 22858 6898
rect 18045 6840 18050 6896
rect 18106 6840 22858 6896
rect 18045 6838 22858 6840
rect 18045 6835 18111 6838
rect 22058 6808 22858 6838
rect 4378 6560 4698 6561
rect 4378 6496 4386 6560
rect 4450 6496 4466 6560
rect 4530 6496 4546 6560
rect 4610 6496 4626 6560
rect 4690 6496 4698 6560
rect 4378 6495 4698 6496
rect 11248 6560 11568 6561
rect 11248 6496 11256 6560
rect 11320 6496 11336 6560
rect 11400 6496 11416 6560
rect 11480 6496 11496 6560
rect 11560 6496 11568 6560
rect 11248 6495 11568 6496
rect 18117 6560 18437 6561
rect 18117 6496 18125 6560
rect 18189 6496 18205 6560
rect 18269 6496 18285 6560
rect 18349 6496 18365 6560
rect 18429 6496 18437 6560
rect 18117 6495 18437 6496
rect 7813 6016 8133 6017
rect 7813 5952 7821 6016
rect 7885 5952 7901 6016
rect 7965 5952 7981 6016
rect 8045 5952 8061 6016
rect 8125 5952 8133 6016
rect 7813 5951 8133 5952
rect 14682 6016 15002 6017
rect 14682 5952 14690 6016
rect 14754 5952 14770 6016
rect 14834 5952 14850 6016
rect 14914 5952 14930 6016
rect 14994 5952 15002 6016
rect 14682 5951 15002 5952
rect 4378 5472 4698 5473
rect 4378 5408 4386 5472
rect 4450 5408 4466 5472
rect 4530 5408 4546 5472
rect 4610 5408 4626 5472
rect 4690 5408 4698 5472
rect 4378 5407 4698 5408
rect 11248 5472 11568 5473
rect 11248 5408 11256 5472
rect 11320 5408 11336 5472
rect 11400 5408 11416 5472
rect 11480 5408 11496 5472
rect 11560 5408 11568 5472
rect 11248 5407 11568 5408
rect 18117 5472 18437 5473
rect 18117 5408 18125 5472
rect 18189 5408 18205 5472
rect 18269 5408 18285 5472
rect 18349 5408 18365 5472
rect 18429 5408 18437 5472
rect 18117 5407 18437 5408
rect 7813 4928 8133 4929
rect 7813 4864 7821 4928
rect 7885 4864 7901 4928
rect 7965 4864 7981 4928
rect 8045 4864 8061 4928
rect 8125 4864 8133 4928
rect 7813 4863 8133 4864
rect 14682 4928 15002 4929
rect 14682 4864 14690 4928
rect 14754 4864 14770 4928
rect 14834 4864 14850 4928
rect 14914 4864 14930 4928
rect 14994 4864 15002 4928
rect 14682 4863 15002 4864
rect 4378 4384 4698 4385
rect 4378 4320 4386 4384
rect 4450 4320 4466 4384
rect 4530 4320 4546 4384
rect 4610 4320 4626 4384
rect 4690 4320 4698 4384
rect 4378 4319 4698 4320
rect 11248 4384 11568 4385
rect 11248 4320 11256 4384
rect 11320 4320 11336 4384
rect 11400 4320 11416 4384
rect 11480 4320 11496 4384
rect 11560 4320 11568 4384
rect 11248 4319 11568 4320
rect 18117 4384 18437 4385
rect 18117 4320 18125 4384
rect 18189 4320 18205 4384
rect 18269 4320 18285 4384
rect 18349 4320 18365 4384
rect 18429 4320 18437 4384
rect 18117 4319 18437 4320
rect 18781 4178 18847 4181
rect 22058 4178 22858 4208
rect 18781 4176 22858 4178
rect 18781 4120 18786 4176
rect 18842 4120 22858 4176
rect 18781 4118 22858 4120
rect 18781 4115 18847 4118
rect 22058 4088 22858 4118
rect 7813 3840 8133 3841
rect 7813 3776 7821 3840
rect 7885 3776 7901 3840
rect 7965 3776 7981 3840
rect 8045 3776 8061 3840
rect 8125 3776 8133 3840
rect 7813 3775 8133 3776
rect 14682 3840 15002 3841
rect 14682 3776 14690 3840
rect 14754 3776 14770 3840
rect 14834 3776 14850 3840
rect 14914 3776 14930 3840
rect 14994 3776 15002 3840
rect 14682 3775 15002 3776
rect 4378 3296 4698 3297
rect 4378 3232 4386 3296
rect 4450 3232 4466 3296
rect 4530 3232 4546 3296
rect 4610 3232 4626 3296
rect 4690 3232 4698 3296
rect 4378 3231 4698 3232
rect 11248 3296 11568 3297
rect 11248 3232 11256 3296
rect 11320 3232 11336 3296
rect 11400 3232 11416 3296
rect 11480 3232 11496 3296
rect 11560 3232 11568 3296
rect 11248 3231 11568 3232
rect 18117 3296 18437 3297
rect 18117 3232 18125 3296
rect 18189 3232 18205 3296
rect 18269 3232 18285 3296
rect 18349 3232 18365 3296
rect 18429 3232 18437 3296
rect 18117 3231 18437 3232
rect 7813 2752 8133 2753
rect 7813 2688 7821 2752
rect 7885 2688 7901 2752
rect 7965 2688 7981 2752
rect 8045 2688 8061 2752
rect 8125 2688 8133 2752
rect 7813 2687 8133 2688
rect 14682 2752 15002 2753
rect 14682 2688 14690 2752
rect 14754 2688 14770 2752
rect 14834 2688 14850 2752
rect 14914 2688 14930 2752
rect 14994 2688 15002 2752
rect 14682 2687 15002 2688
rect 4378 2208 4698 2209
rect 4378 2144 4386 2208
rect 4450 2144 4466 2208
rect 4530 2144 4546 2208
rect 4610 2144 4626 2208
rect 4690 2144 4698 2208
rect 4378 2143 4698 2144
rect 11248 2208 11568 2209
rect 11248 2144 11256 2208
rect 11320 2144 11336 2208
rect 11400 2144 11416 2208
rect 11480 2144 11496 2208
rect 11560 2144 11568 2208
rect 11248 2143 11568 2144
rect 18117 2208 18437 2209
rect 18117 2144 18125 2208
rect 18189 2144 18205 2208
rect 18269 2144 18285 2208
rect 18349 2144 18365 2208
rect 18429 2144 18437 2208
rect 18117 2143 18437 2144
rect 19241 1458 19307 1461
rect 22058 1458 22858 1488
rect 19241 1456 22858 1458
rect 19241 1400 19246 1456
rect 19302 1400 22858 1456
rect 19241 1398 22858 1400
rect 19241 1395 19307 1398
rect 22058 1368 22858 1398
<< via3 >>
rect 7821 22332 7885 22336
rect 7821 22276 7825 22332
rect 7825 22276 7881 22332
rect 7881 22276 7885 22332
rect 7821 22272 7885 22276
rect 7901 22332 7965 22336
rect 7901 22276 7905 22332
rect 7905 22276 7961 22332
rect 7961 22276 7965 22332
rect 7901 22272 7965 22276
rect 7981 22332 8045 22336
rect 7981 22276 7985 22332
rect 7985 22276 8041 22332
rect 8041 22276 8045 22332
rect 7981 22272 8045 22276
rect 8061 22332 8125 22336
rect 8061 22276 8065 22332
rect 8065 22276 8121 22332
rect 8121 22276 8125 22332
rect 8061 22272 8125 22276
rect 14690 22332 14754 22336
rect 14690 22276 14694 22332
rect 14694 22276 14750 22332
rect 14750 22276 14754 22332
rect 14690 22272 14754 22276
rect 14770 22332 14834 22336
rect 14770 22276 14774 22332
rect 14774 22276 14830 22332
rect 14830 22276 14834 22332
rect 14770 22272 14834 22276
rect 14850 22332 14914 22336
rect 14850 22276 14854 22332
rect 14854 22276 14910 22332
rect 14910 22276 14914 22332
rect 14850 22272 14914 22276
rect 14930 22332 14994 22336
rect 14930 22276 14934 22332
rect 14934 22276 14990 22332
rect 14990 22276 14994 22332
rect 14930 22272 14994 22276
rect 4386 21788 4450 21792
rect 4386 21732 4390 21788
rect 4390 21732 4446 21788
rect 4446 21732 4450 21788
rect 4386 21728 4450 21732
rect 4466 21788 4530 21792
rect 4466 21732 4470 21788
rect 4470 21732 4526 21788
rect 4526 21732 4530 21788
rect 4466 21728 4530 21732
rect 4546 21788 4610 21792
rect 4546 21732 4550 21788
rect 4550 21732 4606 21788
rect 4606 21732 4610 21788
rect 4546 21728 4610 21732
rect 4626 21788 4690 21792
rect 4626 21732 4630 21788
rect 4630 21732 4686 21788
rect 4686 21732 4690 21788
rect 4626 21728 4690 21732
rect 11256 21788 11320 21792
rect 11256 21732 11260 21788
rect 11260 21732 11316 21788
rect 11316 21732 11320 21788
rect 11256 21728 11320 21732
rect 11336 21788 11400 21792
rect 11336 21732 11340 21788
rect 11340 21732 11396 21788
rect 11396 21732 11400 21788
rect 11336 21728 11400 21732
rect 11416 21788 11480 21792
rect 11416 21732 11420 21788
rect 11420 21732 11476 21788
rect 11476 21732 11480 21788
rect 11416 21728 11480 21732
rect 11496 21788 11560 21792
rect 11496 21732 11500 21788
rect 11500 21732 11556 21788
rect 11556 21732 11560 21788
rect 11496 21728 11560 21732
rect 18125 21788 18189 21792
rect 18125 21732 18129 21788
rect 18129 21732 18185 21788
rect 18185 21732 18189 21788
rect 18125 21728 18189 21732
rect 18205 21788 18269 21792
rect 18205 21732 18209 21788
rect 18209 21732 18265 21788
rect 18265 21732 18269 21788
rect 18205 21728 18269 21732
rect 18285 21788 18349 21792
rect 18285 21732 18289 21788
rect 18289 21732 18345 21788
rect 18345 21732 18349 21788
rect 18285 21728 18349 21732
rect 18365 21788 18429 21792
rect 18365 21732 18369 21788
rect 18369 21732 18425 21788
rect 18425 21732 18429 21788
rect 18365 21728 18429 21732
rect 7821 21244 7885 21248
rect 7821 21188 7825 21244
rect 7825 21188 7881 21244
rect 7881 21188 7885 21244
rect 7821 21184 7885 21188
rect 7901 21244 7965 21248
rect 7901 21188 7905 21244
rect 7905 21188 7961 21244
rect 7961 21188 7965 21244
rect 7901 21184 7965 21188
rect 7981 21244 8045 21248
rect 7981 21188 7985 21244
rect 7985 21188 8041 21244
rect 8041 21188 8045 21244
rect 7981 21184 8045 21188
rect 8061 21244 8125 21248
rect 8061 21188 8065 21244
rect 8065 21188 8121 21244
rect 8121 21188 8125 21244
rect 8061 21184 8125 21188
rect 14690 21244 14754 21248
rect 14690 21188 14694 21244
rect 14694 21188 14750 21244
rect 14750 21188 14754 21244
rect 14690 21184 14754 21188
rect 14770 21244 14834 21248
rect 14770 21188 14774 21244
rect 14774 21188 14830 21244
rect 14830 21188 14834 21244
rect 14770 21184 14834 21188
rect 14850 21244 14914 21248
rect 14850 21188 14854 21244
rect 14854 21188 14910 21244
rect 14910 21188 14914 21244
rect 14850 21184 14914 21188
rect 14930 21244 14994 21248
rect 14930 21188 14934 21244
rect 14934 21188 14990 21244
rect 14990 21188 14994 21244
rect 14930 21184 14994 21188
rect 4386 20700 4450 20704
rect 4386 20644 4390 20700
rect 4390 20644 4446 20700
rect 4446 20644 4450 20700
rect 4386 20640 4450 20644
rect 4466 20700 4530 20704
rect 4466 20644 4470 20700
rect 4470 20644 4526 20700
rect 4526 20644 4530 20700
rect 4466 20640 4530 20644
rect 4546 20700 4610 20704
rect 4546 20644 4550 20700
rect 4550 20644 4606 20700
rect 4606 20644 4610 20700
rect 4546 20640 4610 20644
rect 4626 20700 4690 20704
rect 4626 20644 4630 20700
rect 4630 20644 4686 20700
rect 4686 20644 4690 20700
rect 4626 20640 4690 20644
rect 11256 20700 11320 20704
rect 11256 20644 11260 20700
rect 11260 20644 11316 20700
rect 11316 20644 11320 20700
rect 11256 20640 11320 20644
rect 11336 20700 11400 20704
rect 11336 20644 11340 20700
rect 11340 20644 11396 20700
rect 11396 20644 11400 20700
rect 11336 20640 11400 20644
rect 11416 20700 11480 20704
rect 11416 20644 11420 20700
rect 11420 20644 11476 20700
rect 11476 20644 11480 20700
rect 11416 20640 11480 20644
rect 11496 20700 11560 20704
rect 11496 20644 11500 20700
rect 11500 20644 11556 20700
rect 11556 20644 11560 20700
rect 11496 20640 11560 20644
rect 18125 20700 18189 20704
rect 18125 20644 18129 20700
rect 18129 20644 18185 20700
rect 18185 20644 18189 20700
rect 18125 20640 18189 20644
rect 18205 20700 18269 20704
rect 18205 20644 18209 20700
rect 18209 20644 18265 20700
rect 18265 20644 18269 20700
rect 18205 20640 18269 20644
rect 18285 20700 18349 20704
rect 18285 20644 18289 20700
rect 18289 20644 18345 20700
rect 18345 20644 18349 20700
rect 18285 20640 18349 20644
rect 18365 20700 18429 20704
rect 18365 20644 18369 20700
rect 18369 20644 18425 20700
rect 18425 20644 18429 20700
rect 18365 20640 18429 20644
rect 7821 20156 7885 20160
rect 7821 20100 7825 20156
rect 7825 20100 7881 20156
rect 7881 20100 7885 20156
rect 7821 20096 7885 20100
rect 7901 20156 7965 20160
rect 7901 20100 7905 20156
rect 7905 20100 7961 20156
rect 7961 20100 7965 20156
rect 7901 20096 7965 20100
rect 7981 20156 8045 20160
rect 7981 20100 7985 20156
rect 7985 20100 8041 20156
rect 8041 20100 8045 20156
rect 7981 20096 8045 20100
rect 8061 20156 8125 20160
rect 8061 20100 8065 20156
rect 8065 20100 8121 20156
rect 8121 20100 8125 20156
rect 8061 20096 8125 20100
rect 14690 20156 14754 20160
rect 14690 20100 14694 20156
rect 14694 20100 14750 20156
rect 14750 20100 14754 20156
rect 14690 20096 14754 20100
rect 14770 20156 14834 20160
rect 14770 20100 14774 20156
rect 14774 20100 14830 20156
rect 14830 20100 14834 20156
rect 14770 20096 14834 20100
rect 14850 20156 14914 20160
rect 14850 20100 14854 20156
rect 14854 20100 14910 20156
rect 14910 20100 14914 20156
rect 14850 20096 14914 20100
rect 14930 20156 14994 20160
rect 14930 20100 14934 20156
rect 14934 20100 14990 20156
rect 14990 20100 14994 20156
rect 14930 20096 14994 20100
rect 4386 19612 4450 19616
rect 4386 19556 4390 19612
rect 4390 19556 4446 19612
rect 4446 19556 4450 19612
rect 4386 19552 4450 19556
rect 4466 19612 4530 19616
rect 4466 19556 4470 19612
rect 4470 19556 4526 19612
rect 4526 19556 4530 19612
rect 4466 19552 4530 19556
rect 4546 19612 4610 19616
rect 4546 19556 4550 19612
rect 4550 19556 4606 19612
rect 4606 19556 4610 19612
rect 4546 19552 4610 19556
rect 4626 19612 4690 19616
rect 4626 19556 4630 19612
rect 4630 19556 4686 19612
rect 4686 19556 4690 19612
rect 4626 19552 4690 19556
rect 11256 19612 11320 19616
rect 11256 19556 11260 19612
rect 11260 19556 11316 19612
rect 11316 19556 11320 19612
rect 11256 19552 11320 19556
rect 11336 19612 11400 19616
rect 11336 19556 11340 19612
rect 11340 19556 11396 19612
rect 11396 19556 11400 19612
rect 11336 19552 11400 19556
rect 11416 19612 11480 19616
rect 11416 19556 11420 19612
rect 11420 19556 11476 19612
rect 11476 19556 11480 19612
rect 11416 19552 11480 19556
rect 11496 19612 11560 19616
rect 11496 19556 11500 19612
rect 11500 19556 11556 19612
rect 11556 19556 11560 19612
rect 11496 19552 11560 19556
rect 18125 19612 18189 19616
rect 18125 19556 18129 19612
rect 18129 19556 18185 19612
rect 18185 19556 18189 19612
rect 18125 19552 18189 19556
rect 18205 19612 18269 19616
rect 18205 19556 18209 19612
rect 18209 19556 18265 19612
rect 18265 19556 18269 19612
rect 18205 19552 18269 19556
rect 18285 19612 18349 19616
rect 18285 19556 18289 19612
rect 18289 19556 18345 19612
rect 18345 19556 18349 19612
rect 18285 19552 18349 19556
rect 18365 19612 18429 19616
rect 18365 19556 18369 19612
rect 18369 19556 18425 19612
rect 18425 19556 18429 19612
rect 18365 19552 18429 19556
rect 7821 19068 7885 19072
rect 7821 19012 7825 19068
rect 7825 19012 7881 19068
rect 7881 19012 7885 19068
rect 7821 19008 7885 19012
rect 7901 19068 7965 19072
rect 7901 19012 7905 19068
rect 7905 19012 7961 19068
rect 7961 19012 7965 19068
rect 7901 19008 7965 19012
rect 7981 19068 8045 19072
rect 7981 19012 7985 19068
rect 7985 19012 8041 19068
rect 8041 19012 8045 19068
rect 7981 19008 8045 19012
rect 8061 19068 8125 19072
rect 8061 19012 8065 19068
rect 8065 19012 8121 19068
rect 8121 19012 8125 19068
rect 8061 19008 8125 19012
rect 14690 19068 14754 19072
rect 14690 19012 14694 19068
rect 14694 19012 14750 19068
rect 14750 19012 14754 19068
rect 14690 19008 14754 19012
rect 14770 19068 14834 19072
rect 14770 19012 14774 19068
rect 14774 19012 14830 19068
rect 14830 19012 14834 19068
rect 14770 19008 14834 19012
rect 14850 19068 14914 19072
rect 14850 19012 14854 19068
rect 14854 19012 14910 19068
rect 14910 19012 14914 19068
rect 14850 19008 14914 19012
rect 14930 19068 14994 19072
rect 14930 19012 14934 19068
rect 14934 19012 14990 19068
rect 14990 19012 14994 19068
rect 14930 19008 14994 19012
rect 4386 18524 4450 18528
rect 4386 18468 4390 18524
rect 4390 18468 4446 18524
rect 4446 18468 4450 18524
rect 4386 18464 4450 18468
rect 4466 18524 4530 18528
rect 4466 18468 4470 18524
rect 4470 18468 4526 18524
rect 4526 18468 4530 18524
rect 4466 18464 4530 18468
rect 4546 18524 4610 18528
rect 4546 18468 4550 18524
rect 4550 18468 4606 18524
rect 4606 18468 4610 18524
rect 4546 18464 4610 18468
rect 4626 18524 4690 18528
rect 4626 18468 4630 18524
rect 4630 18468 4686 18524
rect 4686 18468 4690 18524
rect 4626 18464 4690 18468
rect 11256 18524 11320 18528
rect 11256 18468 11260 18524
rect 11260 18468 11316 18524
rect 11316 18468 11320 18524
rect 11256 18464 11320 18468
rect 11336 18524 11400 18528
rect 11336 18468 11340 18524
rect 11340 18468 11396 18524
rect 11396 18468 11400 18524
rect 11336 18464 11400 18468
rect 11416 18524 11480 18528
rect 11416 18468 11420 18524
rect 11420 18468 11476 18524
rect 11476 18468 11480 18524
rect 11416 18464 11480 18468
rect 11496 18524 11560 18528
rect 11496 18468 11500 18524
rect 11500 18468 11556 18524
rect 11556 18468 11560 18524
rect 11496 18464 11560 18468
rect 18125 18524 18189 18528
rect 18125 18468 18129 18524
rect 18129 18468 18185 18524
rect 18185 18468 18189 18524
rect 18125 18464 18189 18468
rect 18205 18524 18269 18528
rect 18205 18468 18209 18524
rect 18209 18468 18265 18524
rect 18265 18468 18269 18524
rect 18205 18464 18269 18468
rect 18285 18524 18349 18528
rect 18285 18468 18289 18524
rect 18289 18468 18345 18524
rect 18345 18468 18349 18524
rect 18285 18464 18349 18468
rect 18365 18524 18429 18528
rect 18365 18468 18369 18524
rect 18369 18468 18425 18524
rect 18425 18468 18429 18524
rect 18365 18464 18429 18468
rect 7821 17980 7885 17984
rect 7821 17924 7825 17980
rect 7825 17924 7881 17980
rect 7881 17924 7885 17980
rect 7821 17920 7885 17924
rect 7901 17980 7965 17984
rect 7901 17924 7905 17980
rect 7905 17924 7961 17980
rect 7961 17924 7965 17980
rect 7901 17920 7965 17924
rect 7981 17980 8045 17984
rect 7981 17924 7985 17980
rect 7985 17924 8041 17980
rect 8041 17924 8045 17980
rect 7981 17920 8045 17924
rect 8061 17980 8125 17984
rect 8061 17924 8065 17980
rect 8065 17924 8121 17980
rect 8121 17924 8125 17980
rect 8061 17920 8125 17924
rect 14690 17980 14754 17984
rect 14690 17924 14694 17980
rect 14694 17924 14750 17980
rect 14750 17924 14754 17980
rect 14690 17920 14754 17924
rect 14770 17980 14834 17984
rect 14770 17924 14774 17980
rect 14774 17924 14830 17980
rect 14830 17924 14834 17980
rect 14770 17920 14834 17924
rect 14850 17980 14914 17984
rect 14850 17924 14854 17980
rect 14854 17924 14910 17980
rect 14910 17924 14914 17980
rect 14850 17920 14914 17924
rect 14930 17980 14994 17984
rect 14930 17924 14934 17980
rect 14934 17924 14990 17980
rect 14990 17924 14994 17980
rect 14930 17920 14994 17924
rect 4386 17436 4450 17440
rect 4386 17380 4390 17436
rect 4390 17380 4446 17436
rect 4446 17380 4450 17436
rect 4386 17376 4450 17380
rect 4466 17436 4530 17440
rect 4466 17380 4470 17436
rect 4470 17380 4526 17436
rect 4526 17380 4530 17436
rect 4466 17376 4530 17380
rect 4546 17436 4610 17440
rect 4546 17380 4550 17436
rect 4550 17380 4606 17436
rect 4606 17380 4610 17436
rect 4546 17376 4610 17380
rect 4626 17436 4690 17440
rect 4626 17380 4630 17436
rect 4630 17380 4686 17436
rect 4686 17380 4690 17436
rect 4626 17376 4690 17380
rect 11256 17436 11320 17440
rect 11256 17380 11260 17436
rect 11260 17380 11316 17436
rect 11316 17380 11320 17436
rect 11256 17376 11320 17380
rect 11336 17436 11400 17440
rect 11336 17380 11340 17436
rect 11340 17380 11396 17436
rect 11396 17380 11400 17436
rect 11336 17376 11400 17380
rect 11416 17436 11480 17440
rect 11416 17380 11420 17436
rect 11420 17380 11476 17436
rect 11476 17380 11480 17436
rect 11416 17376 11480 17380
rect 11496 17436 11560 17440
rect 11496 17380 11500 17436
rect 11500 17380 11556 17436
rect 11556 17380 11560 17436
rect 11496 17376 11560 17380
rect 18125 17436 18189 17440
rect 18125 17380 18129 17436
rect 18129 17380 18185 17436
rect 18185 17380 18189 17436
rect 18125 17376 18189 17380
rect 18205 17436 18269 17440
rect 18205 17380 18209 17436
rect 18209 17380 18265 17436
rect 18265 17380 18269 17436
rect 18205 17376 18269 17380
rect 18285 17436 18349 17440
rect 18285 17380 18289 17436
rect 18289 17380 18345 17436
rect 18345 17380 18349 17436
rect 18285 17376 18349 17380
rect 18365 17436 18429 17440
rect 18365 17380 18369 17436
rect 18369 17380 18425 17436
rect 18425 17380 18429 17436
rect 18365 17376 18429 17380
rect 7821 16892 7885 16896
rect 7821 16836 7825 16892
rect 7825 16836 7881 16892
rect 7881 16836 7885 16892
rect 7821 16832 7885 16836
rect 7901 16892 7965 16896
rect 7901 16836 7905 16892
rect 7905 16836 7961 16892
rect 7961 16836 7965 16892
rect 7901 16832 7965 16836
rect 7981 16892 8045 16896
rect 7981 16836 7985 16892
rect 7985 16836 8041 16892
rect 8041 16836 8045 16892
rect 7981 16832 8045 16836
rect 8061 16892 8125 16896
rect 8061 16836 8065 16892
rect 8065 16836 8121 16892
rect 8121 16836 8125 16892
rect 8061 16832 8125 16836
rect 14690 16892 14754 16896
rect 14690 16836 14694 16892
rect 14694 16836 14750 16892
rect 14750 16836 14754 16892
rect 14690 16832 14754 16836
rect 14770 16892 14834 16896
rect 14770 16836 14774 16892
rect 14774 16836 14830 16892
rect 14830 16836 14834 16892
rect 14770 16832 14834 16836
rect 14850 16892 14914 16896
rect 14850 16836 14854 16892
rect 14854 16836 14910 16892
rect 14910 16836 14914 16892
rect 14850 16832 14914 16836
rect 14930 16892 14994 16896
rect 14930 16836 14934 16892
rect 14934 16836 14990 16892
rect 14990 16836 14994 16892
rect 14930 16832 14994 16836
rect 4386 16348 4450 16352
rect 4386 16292 4390 16348
rect 4390 16292 4446 16348
rect 4446 16292 4450 16348
rect 4386 16288 4450 16292
rect 4466 16348 4530 16352
rect 4466 16292 4470 16348
rect 4470 16292 4526 16348
rect 4526 16292 4530 16348
rect 4466 16288 4530 16292
rect 4546 16348 4610 16352
rect 4546 16292 4550 16348
rect 4550 16292 4606 16348
rect 4606 16292 4610 16348
rect 4546 16288 4610 16292
rect 4626 16348 4690 16352
rect 4626 16292 4630 16348
rect 4630 16292 4686 16348
rect 4686 16292 4690 16348
rect 4626 16288 4690 16292
rect 11256 16348 11320 16352
rect 11256 16292 11260 16348
rect 11260 16292 11316 16348
rect 11316 16292 11320 16348
rect 11256 16288 11320 16292
rect 11336 16348 11400 16352
rect 11336 16292 11340 16348
rect 11340 16292 11396 16348
rect 11396 16292 11400 16348
rect 11336 16288 11400 16292
rect 11416 16348 11480 16352
rect 11416 16292 11420 16348
rect 11420 16292 11476 16348
rect 11476 16292 11480 16348
rect 11416 16288 11480 16292
rect 11496 16348 11560 16352
rect 11496 16292 11500 16348
rect 11500 16292 11556 16348
rect 11556 16292 11560 16348
rect 11496 16288 11560 16292
rect 18125 16348 18189 16352
rect 18125 16292 18129 16348
rect 18129 16292 18185 16348
rect 18185 16292 18189 16348
rect 18125 16288 18189 16292
rect 18205 16348 18269 16352
rect 18205 16292 18209 16348
rect 18209 16292 18265 16348
rect 18265 16292 18269 16348
rect 18205 16288 18269 16292
rect 18285 16348 18349 16352
rect 18285 16292 18289 16348
rect 18289 16292 18345 16348
rect 18345 16292 18349 16348
rect 18285 16288 18349 16292
rect 18365 16348 18429 16352
rect 18365 16292 18369 16348
rect 18369 16292 18425 16348
rect 18425 16292 18429 16348
rect 18365 16288 18429 16292
rect 7821 15804 7885 15808
rect 7821 15748 7825 15804
rect 7825 15748 7881 15804
rect 7881 15748 7885 15804
rect 7821 15744 7885 15748
rect 7901 15804 7965 15808
rect 7901 15748 7905 15804
rect 7905 15748 7961 15804
rect 7961 15748 7965 15804
rect 7901 15744 7965 15748
rect 7981 15804 8045 15808
rect 7981 15748 7985 15804
rect 7985 15748 8041 15804
rect 8041 15748 8045 15804
rect 7981 15744 8045 15748
rect 8061 15804 8125 15808
rect 8061 15748 8065 15804
rect 8065 15748 8121 15804
rect 8121 15748 8125 15804
rect 8061 15744 8125 15748
rect 14690 15804 14754 15808
rect 14690 15748 14694 15804
rect 14694 15748 14750 15804
rect 14750 15748 14754 15804
rect 14690 15744 14754 15748
rect 14770 15804 14834 15808
rect 14770 15748 14774 15804
rect 14774 15748 14830 15804
rect 14830 15748 14834 15804
rect 14770 15744 14834 15748
rect 14850 15804 14914 15808
rect 14850 15748 14854 15804
rect 14854 15748 14910 15804
rect 14910 15748 14914 15804
rect 14850 15744 14914 15748
rect 14930 15804 14994 15808
rect 14930 15748 14934 15804
rect 14934 15748 14990 15804
rect 14990 15748 14994 15804
rect 14930 15744 14994 15748
rect 4386 15260 4450 15264
rect 4386 15204 4390 15260
rect 4390 15204 4446 15260
rect 4446 15204 4450 15260
rect 4386 15200 4450 15204
rect 4466 15260 4530 15264
rect 4466 15204 4470 15260
rect 4470 15204 4526 15260
rect 4526 15204 4530 15260
rect 4466 15200 4530 15204
rect 4546 15260 4610 15264
rect 4546 15204 4550 15260
rect 4550 15204 4606 15260
rect 4606 15204 4610 15260
rect 4546 15200 4610 15204
rect 4626 15260 4690 15264
rect 4626 15204 4630 15260
rect 4630 15204 4686 15260
rect 4686 15204 4690 15260
rect 4626 15200 4690 15204
rect 11256 15260 11320 15264
rect 11256 15204 11260 15260
rect 11260 15204 11316 15260
rect 11316 15204 11320 15260
rect 11256 15200 11320 15204
rect 11336 15260 11400 15264
rect 11336 15204 11340 15260
rect 11340 15204 11396 15260
rect 11396 15204 11400 15260
rect 11336 15200 11400 15204
rect 11416 15260 11480 15264
rect 11416 15204 11420 15260
rect 11420 15204 11476 15260
rect 11476 15204 11480 15260
rect 11416 15200 11480 15204
rect 11496 15260 11560 15264
rect 11496 15204 11500 15260
rect 11500 15204 11556 15260
rect 11556 15204 11560 15260
rect 11496 15200 11560 15204
rect 18125 15260 18189 15264
rect 18125 15204 18129 15260
rect 18129 15204 18185 15260
rect 18185 15204 18189 15260
rect 18125 15200 18189 15204
rect 18205 15260 18269 15264
rect 18205 15204 18209 15260
rect 18209 15204 18265 15260
rect 18265 15204 18269 15260
rect 18205 15200 18269 15204
rect 18285 15260 18349 15264
rect 18285 15204 18289 15260
rect 18289 15204 18345 15260
rect 18345 15204 18349 15260
rect 18285 15200 18349 15204
rect 18365 15260 18429 15264
rect 18365 15204 18369 15260
rect 18369 15204 18425 15260
rect 18425 15204 18429 15260
rect 18365 15200 18429 15204
rect 7821 14716 7885 14720
rect 7821 14660 7825 14716
rect 7825 14660 7881 14716
rect 7881 14660 7885 14716
rect 7821 14656 7885 14660
rect 7901 14716 7965 14720
rect 7901 14660 7905 14716
rect 7905 14660 7961 14716
rect 7961 14660 7965 14716
rect 7901 14656 7965 14660
rect 7981 14716 8045 14720
rect 7981 14660 7985 14716
rect 7985 14660 8041 14716
rect 8041 14660 8045 14716
rect 7981 14656 8045 14660
rect 8061 14716 8125 14720
rect 8061 14660 8065 14716
rect 8065 14660 8121 14716
rect 8121 14660 8125 14716
rect 8061 14656 8125 14660
rect 14690 14716 14754 14720
rect 14690 14660 14694 14716
rect 14694 14660 14750 14716
rect 14750 14660 14754 14716
rect 14690 14656 14754 14660
rect 14770 14716 14834 14720
rect 14770 14660 14774 14716
rect 14774 14660 14830 14716
rect 14830 14660 14834 14716
rect 14770 14656 14834 14660
rect 14850 14716 14914 14720
rect 14850 14660 14854 14716
rect 14854 14660 14910 14716
rect 14910 14660 14914 14716
rect 14850 14656 14914 14660
rect 14930 14716 14994 14720
rect 14930 14660 14934 14716
rect 14934 14660 14990 14716
rect 14990 14660 14994 14716
rect 14930 14656 14994 14660
rect 4386 14172 4450 14176
rect 4386 14116 4390 14172
rect 4390 14116 4446 14172
rect 4446 14116 4450 14172
rect 4386 14112 4450 14116
rect 4466 14172 4530 14176
rect 4466 14116 4470 14172
rect 4470 14116 4526 14172
rect 4526 14116 4530 14172
rect 4466 14112 4530 14116
rect 4546 14172 4610 14176
rect 4546 14116 4550 14172
rect 4550 14116 4606 14172
rect 4606 14116 4610 14172
rect 4546 14112 4610 14116
rect 4626 14172 4690 14176
rect 4626 14116 4630 14172
rect 4630 14116 4686 14172
rect 4686 14116 4690 14172
rect 4626 14112 4690 14116
rect 11256 14172 11320 14176
rect 11256 14116 11260 14172
rect 11260 14116 11316 14172
rect 11316 14116 11320 14172
rect 11256 14112 11320 14116
rect 11336 14172 11400 14176
rect 11336 14116 11340 14172
rect 11340 14116 11396 14172
rect 11396 14116 11400 14172
rect 11336 14112 11400 14116
rect 11416 14172 11480 14176
rect 11416 14116 11420 14172
rect 11420 14116 11476 14172
rect 11476 14116 11480 14172
rect 11416 14112 11480 14116
rect 11496 14172 11560 14176
rect 11496 14116 11500 14172
rect 11500 14116 11556 14172
rect 11556 14116 11560 14172
rect 11496 14112 11560 14116
rect 18125 14172 18189 14176
rect 18125 14116 18129 14172
rect 18129 14116 18185 14172
rect 18185 14116 18189 14172
rect 18125 14112 18189 14116
rect 18205 14172 18269 14176
rect 18205 14116 18209 14172
rect 18209 14116 18265 14172
rect 18265 14116 18269 14172
rect 18205 14112 18269 14116
rect 18285 14172 18349 14176
rect 18285 14116 18289 14172
rect 18289 14116 18345 14172
rect 18345 14116 18349 14172
rect 18285 14112 18349 14116
rect 18365 14172 18429 14176
rect 18365 14116 18369 14172
rect 18369 14116 18425 14172
rect 18425 14116 18429 14172
rect 18365 14112 18429 14116
rect 7821 13628 7885 13632
rect 7821 13572 7825 13628
rect 7825 13572 7881 13628
rect 7881 13572 7885 13628
rect 7821 13568 7885 13572
rect 7901 13628 7965 13632
rect 7901 13572 7905 13628
rect 7905 13572 7961 13628
rect 7961 13572 7965 13628
rect 7901 13568 7965 13572
rect 7981 13628 8045 13632
rect 7981 13572 7985 13628
rect 7985 13572 8041 13628
rect 8041 13572 8045 13628
rect 7981 13568 8045 13572
rect 8061 13628 8125 13632
rect 8061 13572 8065 13628
rect 8065 13572 8121 13628
rect 8121 13572 8125 13628
rect 8061 13568 8125 13572
rect 14690 13628 14754 13632
rect 14690 13572 14694 13628
rect 14694 13572 14750 13628
rect 14750 13572 14754 13628
rect 14690 13568 14754 13572
rect 14770 13628 14834 13632
rect 14770 13572 14774 13628
rect 14774 13572 14830 13628
rect 14830 13572 14834 13628
rect 14770 13568 14834 13572
rect 14850 13628 14914 13632
rect 14850 13572 14854 13628
rect 14854 13572 14910 13628
rect 14910 13572 14914 13628
rect 14850 13568 14914 13572
rect 14930 13628 14994 13632
rect 14930 13572 14934 13628
rect 14934 13572 14990 13628
rect 14990 13572 14994 13628
rect 14930 13568 14994 13572
rect 4386 13084 4450 13088
rect 4386 13028 4390 13084
rect 4390 13028 4446 13084
rect 4446 13028 4450 13084
rect 4386 13024 4450 13028
rect 4466 13084 4530 13088
rect 4466 13028 4470 13084
rect 4470 13028 4526 13084
rect 4526 13028 4530 13084
rect 4466 13024 4530 13028
rect 4546 13084 4610 13088
rect 4546 13028 4550 13084
rect 4550 13028 4606 13084
rect 4606 13028 4610 13084
rect 4546 13024 4610 13028
rect 4626 13084 4690 13088
rect 4626 13028 4630 13084
rect 4630 13028 4686 13084
rect 4686 13028 4690 13084
rect 4626 13024 4690 13028
rect 11256 13084 11320 13088
rect 11256 13028 11260 13084
rect 11260 13028 11316 13084
rect 11316 13028 11320 13084
rect 11256 13024 11320 13028
rect 11336 13084 11400 13088
rect 11336 13028 11340 13084
rect 11340 13028 11396 13084
rect 11396 13028 11400 13084
rect 11336 13024 11400 13028
rect 11416 13084 11480 13088
rect 11416 13028 11420 13084
rect 11420 13028 11476 13084
rect 11476 13028 11480 13084
rect 11416 13024 11480 13028
rect 11496 13084 11560 13088
rect 11496 13028 11500 13084
rect 11500 13028 11556 13084
rect 11556 13028 11560 13084
rect 11496 13024 11560 13028
rect 18125 13084 18189 13088
rect 18125 13028 18129 13084
rect 18129 13028 18185 13084
rect 18185 13028 18189 13084
rect 18125 13024 18189 13028
rect 18205 13084 18269 13088
rect 18205 13028 18209 13084
rect 18209 13028 18265 13084
rect 18265 13028 18269 13084
rect 18205 13024 18269 13028
rect 18285 13084 18349 13088
rect 18285 13028 18289 13084
rect 18289 13028 18345 13084
rect 18345 13028 18349 13084
rect 18285 13024 18349 13028
rect 18365 13084 18429 13088
rect 18365 13028 18369 13084
rect 18369 13028 18425 13084
rect 18425 13028 18429 13084
rect 18365 13024 18429 13028
rect 7821 12540 7885 12544
rect 7821 12484 7825 12540
rect 7825 12484 7881 12540
rect 7881 12484 7885 12540
rect 7821 12480 7885 12484
rect 7901 12540 7965 12544
rect 7901 12484 7905 12540
rect 7905 12484 7961 12540
rect 7961 12484 7965 12540
rect 7901 12480 7965 12484
rect 7981 12540 8045 12544
rect 7981 12484 7985 12540
rect 7985 12484 8041 12540
rect 8041 12484 8045 12540
rect 7981 12480 8045 12484
rect 8061 12540 8125 12544
rect 8061 12484 8065 12540
rect 8065 12484 8121 12540
rect 8121 12484 8125 12540
rect 8061 12480 8125 12484
rect 14690 12540 14754 12544
rect 14690 12484 14694 12540
rect 14694 12484 14750 12540
rect 14750 12484 14754 12540
rect 14690 12480 14754 12484
rect 14770 12540 14834 12544
rect 14770 12484 14774 12540
rect 14774 12484 14830 12540
rect 14830 12484 14834 12540
rect 14770 12480 14834 12484
rect 14850 12540 14914 12544
rect 14850 12484 14854 12540
rect 14854 12484 14910 12540
rect 14910 12484 14914 12540
rect 14850 12480 14914 12484
rect 14930 12540 14994 12544
rect 14930 12484 14934 12540
rect 14934 12484 14990 12540
rect 14990 12484 14994 12540
rect 14930 12480 14994 12484
rect 4386 11996 4450 12000
rect 4386 11940 4390 11996
rect 4390 11940 4446 11996
rect 4446 11940 4450 11996
rect 4386 11936 4450 11940
rect 4466 11996 4530 12000
rect 4466 11940 4470 11996
rect 4470 11940 4526 11996
rect 4526 11940 4530 11996
rect 4466 11936 4530 11940
rect 4546 11996 4610 12000
rect 4546 11940 4550 11996
rect 4550 11940 4606 11996
rect 4606 11940 4610 11996
rect 4546 11936 4610 11940
rect 4626 11996 4690 12000
rect 4626 11940 4630 11996
rect 4630 11940 4686 11996
rect 4686 11940 4690 11996
rect 4626 11936 4690 11940
rect 11256 11996 11320 12000
rect 11256 11940 11260 11996
rect 11260 11940 11316 11996
rect 11316 11940 11320 11996
rect 11256 11936 11320 11940
rect 11336 11996 11400 12000
rect 11336 11940 11340 11996
rect 11340 11940 11396 11996
rect 11396 11940 11400 11996
rect 11336 11936 11400 11940
rect 11416 11996 11480 12000
rect 11416 11940 11420 11996
rect 11420 11940 11476 11996
rect 11476 11940 11480 11996
rect 11416 11936 11480 11940
rect 11496 11996 11560 12000
rect 11496 11940 11500 11996
rect 11500 11940 11556 11996
rect 11556 11940 11560 11996
rect 11496 11936 11560 11940
rect 18125 11996 18189 12000
rect 18125 11940 18129 11996
rect 18129 11940 18185 11996
rect 18185 11940 18189 11996
rect 18125 11936 18189 11940
rect 18205 11996 18269 12000
rect 18205 11940 18209 11996
rect 18209 11940 18265 11996
rect 18265 11940 18269 11996
rect 18205 11936 18269 11940
rect 18285 11996 18349 12000
rect 18285 11940 18289 11996
rect 18289 11940 18345 11996
rect 18345 11940 18349 11996
rect 18285 11936 18349 11940
rect 18365 11996 18429 12000
rect 18365 11940 18369 11996
rect 18369 11940 18425 11996
rect 18425 11940 18429 11996
rect 18365 11936 18429 11940
rect 7821 11452 7885 11456
rect 7821 11396 7825 11452
rect 7825 11396 7881 11452
rect 7881 11396 7885 11452
rect 7821 11392 7885 11396
rect 7901 11452 7965 11456
rect 7901 11396 7905 11452
rect 7905 11396 7961 11452
rect 7961 11396 7965 11452
rect 7901 11392 7965 11396
rect 7981 11452 8045 11456
rect 7981 11396 7985 11452
rect 7985 11396 8041 11452
rect 8041 11396 8045 11452
rect 7981 11392 8045 11396
rect 8061 11452 8125 11456
rect 8061 11396 8065 11452
rect 8065 11396 8121 11452
rect 8121 11396 8125 11452
rect 8061 11392 8125 11396
rect 14690 11452 14754 11456
rect 14690 11396 14694 11452
rect 14694 11396 14750 11452
rect 14750 11396 14754 11452
rect 14690 11392 14754 11396
rect 14770 11452 14834 11456
rect 14770 11396 14774 11452
rect 14774 11396 14830 11452
rect 14830 11396 14834 11452
rect 14770 11392 14834 11396
rect 14850 11452 14914 11456
rect 14850 11396 14854 11452
rect 14854 11396 14910 11452
rect 14910 11396 14914 11452
rect 14850 11392 14914 11396
rect 14930 11452 14994 11456
rect 14930 11396 14934 11452
rect 14934 11396 14990 11452
rect 14990 11396 14994 11452
rect 14930 11392 14994 11396
rect 4386 10908 4450 10912
rect 4386 10852 4390 10908
rect 4390 10852 4446 10908
rect 4446 10852 4450 10908
rect 4386 10848 4450 10852
rect 4466 10908 4530 10912
rect 4466 10852 4470 10908
rect 4470 10852 4526 10908
rect 4526 10852 4530 10908
rect 4466 10848 4530 10852
rect 4546 10908 4610 10912
rect 4546 10852 4550 10908
rect 4550 10852 4606 10908
rect 4606 10852 4610 10908
rect 4546 10848 4610 10852
rect 4626 10908 4690 10912
rect 4626 10852 4630 10908
rect 4630 10852 4686 10908
rect 4686 10852 4690 10908
rect 4626 10848 4690 10852
rect 11256 10908 11320 10912
rect 11256 10852 11260 10908
rect 11260 10852 11316 10908
rect 11316 10852 11320 10908
rect 11256 10848 11320 10852
rect 11336 10908 11400 10912
rect 11336 10852 11340 10908
rect 11340 10852 11396 10908
rect 11396 10852 11400 10908
rect 11336 10848 11400 10852
rect 11416 10908 11480 10912
rect 11416 10852 11420 10908
rect 11420 10852 11476 10908
rect 11476 10852 11480 10908
rect 11416 10848 11480 10852
rect 11496 10908 11560 10912
rect 11496 10852 11500 10908
rect 11500 10852 11556 10908
rect 11556 10852 11560 10908
rect 11496 10848 11560 10852
rect 18125 10908 18189 10912
rect 18125 10852 18129 10908
rect 18129 10852 18185 10908
rect 18185 10852 18189 10908
rect 18125 10848 18189 10852
rect 18205 10908 18269 10912
rect 18205 10852 18209 10908
rect 18209 10852 18265 10908
rect 18265 10852 18269 10908
rect 18205 10848 18269 10852
rect 18285 10908 18349 10912
rect 18285 10852 18289 10908
rect 18289 10852 18345 10908
rect 18345 10852 18349 10908
rect 18285 10848 18349 10852
rect 18365 10908 18429 10912
rect 18365 10852 18369 10908
rect 18369 10852 18425 10908
rect 18425 10852 18429 10908
rect 18365 10848 18429 10852
rect 7821 10364 7885 10368
rect 7821 10308 7825 10364
rect 7825 10308 7881 10364
rect 7881 10308 7885 10364
rect 7821 10304 7885 10308
rect 7901 10364 7965 10368
rect 7901 10308 7905 10364
rect 7905 10308 7961 10364
rect 7961 10308 7965 10364
rect 7901 10304 7965 10308
rect 7981 10364 8045 10368
rect 7981 10308 7985 10364
rect 7985 10308 8041 10364
rect 8041 10308 8045 10364
rect 7981 10304 8045 10308
rect 8061 10364 8125 10368
rect 8061 10308 8065 10364
rect 8065 10308 8121 10364
rect 8121 10308 8125 10364
rect 8061 10304 8125 10308
rect 14690 10364 14754 10368
rect 14690 10308 14694 10364
rect 14694 10308 14750 10364
rect 14750 10308 14754 10364
rect 14690 10304 14754 10308
rect 14770 10364 14834 10368
rect 14770 10308 14774 10364
rect 14774 10308 14830 10364
rect 14830 10308 14834 10364
rect 14770 10304 14834 10308
rect 14850 10364 14914 10368
rect 14850 10308 14854 10364
rect 14854 10308 14910 10364
rect 14910 10308 14914 10364
rect 14850 10304 14914 10308
rect 14930 10364 14994 10368
rect 14930 10308 14934 10364
rect 14934 10308 14990 10364
rect 14990 10308 14994 10364
rect 14930 10304 14994 10308
rect 4386 9820 4450 9824
rect 4386 9764 4390 9820
rect 4390 9764 4446 9820
rect 4446 9764 4450 9820
rect 4386 9760 4450 9764
rect 4466 9820 4530 9824
rect 4466 9764 4470 9820
rect 4470 9764 4526 9820
rect 4526 9764 4530 9820
rect 4466 9760 4530 9764
rect 4546 9820 4610 9824
rect 4546 9764 4550 9820
rect 4550 9764 4606 9820
rect 4606 9764 4610 9820
rect 4546 9760 4610 9764
rect 4626 9820 4690 9824
rect 4626 9764 4630 9820
rect 4630 9764 4686 9820
rect 4686 9764 4690 9820
rect 4626 9760 4690 9764
rect 11256 9820 11320 9824
rect 11256 9764 11260 9820
rect 11260 9764 11316 9820
rect 11316 9764 11320 9820
rect 11256 9760 11320 9764
rect 11336 9820 11400 9824
rect 11336 9764 11340 9820
rect 11340 9764 11396 9820
rect 11396 9764 11400 9820
rect 11336 9760 11400 9764
rect 11416 9820 11480 9824
rect 11416 9764 11420 9820
rect 11420 9764 11476 9820
rect 11476 9764 11480 9820
rect 11416 9760 11480 9764
rect 11496 9820 11560 9824
rect 11496 9764 11500 9820
rect 11500 9764 11556 9820
rect 11556 9764 11560 9820
rect 11496 9760 11560 9764
rect 18125 9820 18189 9824
rect 18125 9764 18129 9820
rect 18129 9764 18185 9820
rect 18185 9764 18189 9820
rect 18125 9760 18189 9764
rect 18205 9820 18269 9824
rect 18205 9764 18209 9820
rect 18209 9764 18265 9820
rect 18265 9764 18269 9820
rect 18205 9760 18269 9764
rect 18285 9820 18349 9824
rect 18285 9764 18289 9820
rect 18289 9764 18345 9820
rect 18345 9764 18349 9820
rect 18285 9760 18349 9764
rect 18365 9820 18429 9824
rect 18365 9764 18369 9820
rect 18369 9764 18425 9820
rect 18425 9764 18429 9820
rect 18365 9760 18429 9764
rect 7821 9276 7885 9280
rect 7821 9220 7825 9276
rect 7825 9220 7881 9276
rect 7881 9220 7885 9276
rect 7821 9216 7885 9220
rect 7901 9276 7965 9280
rect 7901 9220 7905 9276
rect 7905 9220 7961 9276
rect 7961 9220 7965 9276
rect 7901 9216 7965 9220
rect 7981 9276 8045 9280
rect 7981 9220 7985 9276
rect 7985 9220 8041 9276
rect 8041 9220 8045 9276
rect 7981 9216 8045 9220
rect 8061 9276 8125 9280
rect 8061 9220 8065 9276
rect 8065 9220 8121 9276
rect 8121 9220 8125 9276
rect 8061 9216 8125 9220
rect 14690 9276 14754 9280
rect 14690 9220 14694 9276
rect 14694 9220 14750 9276
rect 14750 9220 14754 9276
rect 14690 9216 14754 9220
rect 14770 9276 14834 9280
rect 14770 9220 14774 9276
rect 14774 9220 14830 9276
rect 14830 9220 14834 9276
rect 14770 9216 14834 9220
rect 14850 9276 14914 9280
rect 14850 9220 14854 9276
rect 14854 9220 14910 9276
rect 14910 9220 14914 9276
rect 14850 9216 14914 9220
rect 14930 9276 14994 9280
rect 14930 9220 14934 9276
rect 14934 9220 14990 9276
rect 14990 9220 14994 9276
rect 14930 9216 14994 9220
rect 4386 8732 4450 8736
rect 4386 8676 4390 8732
rect 4390 8676 4446 8732
rect 4446 8676 4450 8732
rect 4386 8672 4450 8676
rect 4466 8732 4530 8736
rect 4466 8676 4470 8732
rect 4470 8676 4526 8732
rect 4526 8676 4530 8732
rect 4466 8672 4530 8676
rect 4546 8732 4610 8736
rect 4546 8676 4550 8732
rect 4550 8676 4606 8732
rect 4606 8676 4610 8732
rect 4546 8672 4610 8676
rect 4626 8732 4690 8736
rect 4626 8676 4630 8732
rect 4630 8676 4686 8732
rect 4686 8676 4690 8732
rect 4626 8672 4690 8676
rect 11256 8732 11320 8736
rect 11256 8676 11260 8732
rect 11260 8676 11316 8732
rect 11316 8676 11320 8732
rect 11256 8672 11320 8676
rect 11336 8732 11400 8736
rect 11336 8676 11340 8732
rect 11340 8676 11396 8732
rect 11396 8676 11400 8732
rect 11336 8672 11400 8676
rect 11416 8732 11480 8736
rect 11416 8676 11420 8732
rect 11420 8676 11476 8732
rect 11476 8676 11480 8732
rect 11416 8672 11480 8676
rect 11496 8732 11560 8736
rect 11496 8676 11500 8732
rect 11500 8676 11556 8732
rect 11556 8676 11560 8732
rect 11496 8672 11560 8676
rect 18125 8732 18189 8736
rect 18125 8676 18129 8732
rect 18129 8676 18185 8732
rect 18185 8676 18189 8732
rect 18125 8672 18189 8676
rect 18205 8732 18269 8736
rect 18205 8676 18209 8732
rect 18209 8676 18265 8732
rect 18265 8676 18269 8732
rect 18205 8672 18269 8676
rect 18285 8732 18349 8736
rect 18285 8676 18289 8732
rect 18289 8676 18345 8732
rect 18345 8676 18349 8732
rect 18285 8672 18349 8676
rect 18365 8732 18429 8736
rect 18365 8676 18369 8732
rect 18369 8676 18425 8732
rect 18425 8676 18429 8732
rect 18365 8672 18429 8676
rect 7821 8188 7885 8192
rect 7821 8132 7825 8188
rect 7825 8132 7881 8188
rect 7881 8132 7885 8188
rect 7821 8128 7885 8132
rect 7901 8188 7965 8192
rect 7901 8132 7905 8188
rect 7905 8132 7961 8188
rect 7961 8132 7965 8188
rect 7901 8128 7965 8132
rect 7981 8188 8045 8192
rect 7981 8132 7985 8188
rect 7985 8132 8041 8188
rect 8041 8132 8045 8188
rect 7981 8128 8045 8132
rect 8061 8188 8125 8192
rect 8061 8132 8065 8188
rect 8065 8132 8121 8188
rect 8121 8132 8125 8188
rect 8061 8128 8125 8132
rect 14690 8188 14754 8192
rect 14690 8132 14694 8188
rect 14694 8132 14750 8188
rect 14750 8132 14754 8188
rect 14690 8128 14754 8132
rect 14770 8188 14834 8192
rect 14770 8132 14774 8188
rect 14774 8132 14830 8188
rect 14830 8132 14834 8188
rect 14770 8128 14834 8132
rect 14850 8188 14914 8192
rect 14850 8132 14854 8188
rect 14854 8132 14910 8188
rect 14910 8132 14914 8188
rect 14850 8128 14914 8132
rect 14930 8188 14994 8192
rect 14930 8132 14934 8188
rect 14934 8132 14990 8188
rect 14990 8132 14994 8188
rect 14930 8128 14994 8132
rect 4386 7644 4450 7648
rect 4386 7588 4390 7644
rect 4390 7588 4446 7644
rect 4446 7588 4450 7644
rect 4386 7584 4450 7588
rect 4466 7644 4530 7648
rect 4466 7588 4470 7644
rect 4470 7588 4526 7644
rect 4526 7588 4530 7644
rect 4466 7584 4530 7588
rect 4546 7644 4610 7648
rect 4546 7588 4550 7644
rect 4550 7588 4606 7644
rect 4606 7588 4610 7644
rect 4546 7584 4610 7588
rect 4626 7644 4690 7648
rect 4626 7588 4630 7644
rect 4630 7588 4686 7644
rect 4686 7588 4690 7644
rect 4626 7584 4690 7588
rect 11256 7644 11320 7648
rect 11256 7588 11260 7644
rect 11260 7588 11316 7644
rect 11316 7588 11320 7644
rect 11256 7584 11320 7588
rect 11336 7644 11400 7648
rect 11336 7588 11340 7644
rect 11340 7588 11396 7644
rect 11396 7588 11400 7644
rect 11336 7584 11400 7588
rect 11416 7644 11480 7648
rect 11416 7588 11420 7644
rect 11420 7588 11476 7644
rect 11476 7588 11480 7644
rect 11416 7584 11480 7588
rect 11496 7644 11560 7648
rect 11496 7588 11500 7644
rect 11500 7588 11556 7644
rect 11556 7588 11560 7644
rect 11496 7584 11560 7588
rect 18125 7644 18189 7648
rect 18125 7588 18129 7644
rect 18129 7588 18185 7644
rect 18185 7588 18189 7644
rect 18125 7584 18189 7588
rect 18205 7644 18269 7648
rect 18205 7588 18209 7644
rect 18209 7588 18265 7644
rect 18265 7588 18269 7644
rect 18205 7584 18269 7588
rect 18285 7644 18349 7648
rect 18285 7588 18289 7644
rect 18289 7588 18345 7644
rect 18345 7588 18349 7644
rect 18285 7584 18349 7588
rect 18365 7644 18429 7648
rect 18365 7588 18369 7644
rect 18369 7588 18425 7644
rect 18425 7588 18429 7644
rect 18365 7584 18429 7588
rect 7821 7100 7885 7104
rect 7821 7044 7825 7100
rect 7825 7044 7881 7100
rect 7881 7044 7885 7100
rect 7821 7040 7885 7044
rect 7901 7100 7965 7104
rect 7901 7044 7905 7100
rect 7905 7044 7961 7100
rect 7961 7044 7965 7100
rect 7901 7040 7965 7044
rect 7981 7100 8045 7104
rect 7981 7044 7985 7100
rect 7985 7044 8041 7100
rect 8041 7044 8045 7100
rect 7981 7040 8045 7044
rect 8061 7100 8125 7104
rect 8061 7044 8065 7100
rect 8065 7044 8121 7100
rect 8121 7044 8125 7100
rect 8061 7040 8125 7044
rect 14690 7100 14754 7104
rect 14690 7044 14694 7100
rect 14694 7044 14750 7100
rect 14750 7044 14754 7100
rect 14690 7040 14754 7044
rect 14770 7100 14834 7104
rect 14770 7044 14774 7100
rect 14774 7044 14830 7100
rect 14830 7044 14834 7100
rect 14770 7040 14834 7044
rect 14850 7100 14914 7104
rect 14850 7044 14854 7100
rect 14854 7044 14910 7100
rect 14910 7044 14914 7100
rect 14850 7040 14914 7044
rect 14930 7100 14994 7104
rect 14930 7044 14934 7100
rect 14934 7044 14990 7100
rect 14990 7044 14994 7100
rect 14930 7040 14994 7044
rect 4386 6556 4450 6560
rect 4386 6500 4390 6556
rect 4390 6500 4446 6556
rect 4446 6500 4450 6556
rect 4386 6496 4450 6500
rect 4466 6556 4530 6560
rect 4466 6500 4470 6556
rect 4470 6500 4526 6556
rect 4526 6500 4530 6556
rect 4466 6496 4530 6500
rect 4546 6556 4610 6560
rect 4546 6500 4550 6556
rect 4550 6500 4606 6556
rect 4606 6500 4610 6556
rect 4546 6496 4610 6500
rect 4626 6556 4690 6560
rect 4626 6500 4630 6556
rect 4630 6500 4686 6556
rect 4686 6500 4690 6556
rect 4626 6496 4690 6500
rect 11256 6556 11320 6560
rect 11256 6500 11260 6556
rect 11260 6500 11316 6556
rect 11316 6500 11320 6556
rect 11256 6496 11320 6500
rect 11336 6556 11400 6560
rect 11336 6500 11340 6556
rect 11340 6500 11396 6556
rect 11396 6500 11400 6556
rect 11336 6496 11400 6500
rect 11416 6556 11480 6560
rect 11416 6500 11420 6556
rect 11420 6500 11476 6556
rect 11476 6500 11480 6556
rect 11416 6496 11480 6500
rect 11496 6556 11560 6560
rect 11496 6500 11500 6556
rect 11500 6500 11556 6556
rect 11556 6500 11560 6556
rect 11496 6496 11560 6500
rect 18125 6556 18189 6560
rect 18125 6500 18129 6556
rect 18129 6500 18185 6556
rect 18185 6500 18189 6556
rect 18125 6496 18189 6500
rect 18205 6556 18269 6560
rect 18205 6500 18209 6556
rect 18209 6500 18265 6556
rect 18265 6500 18269 6556
rect 18205 6496 18269 6500
rect 18285 6556 18349 6560
rect 18285 6500 18289 6556
rect 18289 6500 18345 6556
rect 18345 6500 18349 6556
rect 18285 6496 18349 6500
rect 18365 6556 18429 6560
rect 18365 6500 18369 6556
rect 18369 6500 18425 6556
rect 18425 6500 18429 6556
rect 18365 6496 18429 6500
rect 7821 6012 7885 6016
rect 7821 5956 7825 6012
rect 7825 5956 7881 6012
rect 7881 5956 7885 6012
rect 7821 5952 7885 5956
rect 7901 6012 7965 6016
rect 7901 5956 7905 6012
rect 7905 5956 7961 6012
rect 7961 5956 7965 6012
rect 7901 5952 7965 5956
rect 7981 6012 8045 6016
rect 7981 5956 7985 6012
rect 7985 5956 8041 6012
rect 8041 5956 8045 6012
rect 7981 5952 8045 5956
rect 8061 6012 8125 6016
rect 8061 5956 8065 6012
rect 8065 5956 8121 6012
rect 8121 5956 8125 6012
rect 8061 5952 8125 5956
rect 14690 6012 14754 6016
rect 14690 5956 14694 6012
rect 14694 5956 14750 6012
rect 14750 5956 14754 6012
rect 14690 5952 14754 5956
rect 14770 6012 14834 6016
rect 14770 5956 14774 6012
rect 14774 5956 14830 6012
rect 14830 5956 14834 6012
rect 14770 5952 14834 5956
rect 14850 6012 14914 6016
rect 14850 5956 14854 6012
rect 14854 5956 14910 6012
rect 14910 5956 14914 6012
rect 14850 5952 14914 5956
rect 14930 6012 14994 6016
rect 14930 5956 14934 6012
rect 14934 5956 14990 6012
rect 14990 5956 14994 6012
rect 14930 5952 14994 5956
rect 4386 5468 4450 5472
rect 4386 5412 4390 5468
rect 4390 5412 4446 5468
rect 4446 5412 4450 5468
rect 4386 5408 4450 5412
rect 4466 5468 4530 5472
rect 4466 5412 4470 5468
rect 4470 5412 4526 5468
rect 4526 5412 4530 5468
rect 4466 5408 4530 5412
rect 4546 5468 4610 5472
rect 4546 5412 4550 5468
rect 4550 5412 4606 5468
rect 4606 5412 4610 5468
rect 4546 5408 4610 5412
rect 4626 5468 4690 5472
rect 4626 5412 4630 5468
rect 4630 5412 4686 5468
rect 4686 5412 4690 5468
rect 4626 5408 4690 5412
rect 11256 5468 11320 5472
rect 11256 5412 11260 5468
rect 11260 5412 11316 5468
rect 11316 5412 11320 5468
rect 11256 5408 11320 5412
rect 11336 5468 11400 5472
rect 11336 5412 11340 5468
rect 11340 5412 11396 5468
rect 11396 5412 11400 5468
rect 11336 5408 11400 5412
rect 11416 5468 11480 5472
rect 11416 5412 11420 5468
rect 11420 5412 11476 5468
rect 11476 5412 11480 5468
rect 11416 5408 11480 5412
rect 11496 5468 11560 5472
rect 11496 5412 11500 5468
rect 11500 5412 11556 5468
rect 11556 5412 11560 5468
rect 11496 5408 11560 5412
rect 18125 5468 18189 5472
rect 18125 5412 18129 5468
rect 18129 5412 18185 5468
rect 18185 5412 18189 5468
rect 18125 5408 18189 5412
rect 18205 5468 18269 5472
rect 18205 5412 18209 5468
rect 18209 5412 18265 5468
rect 18265 5412 18269 5468
rect 18205 5408 18269 5412
rect 18285 5468 18349 5472
rect 18285 5412 18289 5468
rect 18289 5412 18345 5468
rect 18345 5412 18349 5468
rect 18285 5408 18349 5412
rect 18365 5468 18429 5472
rect 18365 5412 18369 5468
rect 18369 5412 18425 5468
rect 18425 5412 18429 5468
rect 18365 5408 18429 5412
rect 7821 4924 7885 4928
rect 7821 4868 7825 4924
rect 7825 4868 7881 4924
rect 7881 4868 7885 4924
rect 7821 4864 7885 4868
rect 7901 4924 7965 4928
rect 7901 4868 7905 4924
rect 7905 4868 7961 4924
rect 7961 4868 7965 4924
rect 7901 4864 7965 4868
rect 7981 4924 8045 4928
rect 7981 4868 7985 4924
rect 7985 4868 8041 4924
rect 8041 4868 8045 4924
rect 7981 4864 8045 4868
rect 8061 4924 8125 4928
rect 8061 4868 8065 4924
rect 8065 4868 8121 4924
rect 8121 4868 8125 4924
rect 8061 4864 8125 4868
rect 14690 4924 14754 4928
rect 14690 4868 14694 4924
rect 14694 4868 14750 4924
rect 14750 4868 14754 4924
rect 14690 4864 14754 4868
rect 14770 4924 14834 4928
rect 14770 4868 14774 4924
rect 14774 4868 14830 4924
rect 14830 4868 14834 4924
rect 14770 4864 14834 4868
rect 14850 4924 14914 4928
rect 14850 4868 14854 4924
rect 14854 4868 14910 4924
rect 14910 4868 14914 4924
rect 14850 4864 14914 4868
rect 14930 4924 14994 4928
rect 14930 4868 14934 4924
rect 14934 4868 14990 4924
rect 14990 4868 14994 4924
rect 14930 4864 14994 4868
rect 4386 4380 4450 4384
rect 4386 4324 4390 4380
rect 4390 4324 4446 4380
rect 4446 4324 4450 4380
rect 4386 4320 4450 4324
rect 4466 4380 4530 4384
rect 4466 4324 4470 4380
rect 4470 4324 4526 4380
rect 4526 4324 4530 4380
rect 4466 4320 4530 4324
rect 4546 4380 4610 4384
rect 4546 4324 4550 4380
rect 4550 4324 4606 4380
rect 4606 4324 4610 4380
rect 4546 4320 4610 4324
rect 4626 4380 4690 4384
rect 4626 4324 4630 4380
rect 4630 4324 4686 4380
rect 4686 4324 4690 4380
rect 4626 4320 4690 4324
rect 11256 4380 11320 4384
rect 11256 4324 11260 4380
rect 11260 4324 11316 4380
rect 11316 4324 11320 4380
rect 11256 4320 11320 4324
rect 11336 4380 11400 4384
rect 11336 4324 11340 4380
rect 11340 4324 11396 4380
rect 11396 4324 11400 4380
rect 11336 4320 11400 4324
rect 11416 4380 11480 4384
rect 11416 4324 11420 4380
rect 11420 4324 11476 4380
rect 11476 4324 11480 4380
rect 11416 4320 11480 4324
rect 11496 4380 11560 4384
rect 11496 4324 11500 4380
rect 11500 4324 11556 4380
rect 11556 4324 11560 4380
rect 11496 4320 11560 4324
rect 18125 4380 18189 4384
rect 18125 4324 18129 4380
rect 18129 4324 18185 4380
rect 18185 4324 18189 4380
rect 18125 4320 18189 4324
rect 18205 4380 18269 4384
rect 18205 4324 18209 4380
rect 18209 4324 18265 4380
rect 18265 4324 18269 4380
rect 18205 4320 18269 4324
rect 18285 4380 18349 4384
rect 18285 4324 18289 4380
rect 18289 4324 18345 4380
rect 18345 4324 18349 4380
rect 18285 4320 18349 4324
rect 18365 4380 18429 4384
rect 18365 4324 18369 4380
rect 18369 4324 18425 4380
rect 18425 4324 18429 4380
rect 18365 4320 18429 4324
rect 7821 3836 7885 3840
rect 7821 3780 7825 3836
rect 7825 3780 7881 3836
rect 7881 3780 7885 3836
rect 7821 3776 7885 3780
rect 7901 3836 7965 3840
rect 7901 3780 7905 3836
rect 7905 3780 7961 3836
rect 7961 3780 7965 3836
rect 7901 3776 7965 3780
rect 7981 3836 8045 3840
rect 7981 3780 7985 3836
rect 7985 3780 8041 3836
rect 8041 3780 8045 3836
rect 7981 3776 8045 3780
rect 8061 3836 8125 3840
rect 8061 3780 8065 3836
rect 8065 3780 8121 3836
rect 8121 3780 8125 3836
rect 8061 3776 8125 3780
rect 14690 3836 14754 3840
rect 14690 3780 14694 3836
rect 14694 3780 14750 3836
rect 14750 3780 14754 3836
rect 14690 3776 14754 3780
rect 14770 3836 14834 3840
rect 14770 3780 14774 3836
rect 14774 3780 14830 3836
rect 14830 3780 14834 3836
rect 14770 3776 14834 3780
rect 14850 3836 14914 3840
rect 14850 3780 14854 3836
rect 14854 3780 14910 3836
rect 14910 3780 14914 3836
rect 14850 3776 14914 3780
rect 14930 3836 14994 3840
rect 14930 3780 14934 3836
rect 14934 3780 14990 3836
rect 14990 3780 14994 3836
rect 14930 3776 14994 3780
rect 4386 3292 4450 3296
rect 4386 3236 4390 3292
rect 4390 3236 4446 3292
rect 4446 3236 4450 3292
rect 4386 3232 4450 3236
rect 4466 3292 4530 3296
rect 4466 3236 4470 3292
rect 4470 3236 4526 3292
rect 4526 3236 4530 3292
rect 4466 3232 4530 3236
rect 4546 3292 4610 3296
rect 4546 3236 4550 3292
rect 4550 3236 4606 3292
rect 4606 3236 4610 3292
rect 4546 3232 4610 3236
rect 4626 3292 4690 3296
rect 4626 3236 4630 3292
rect 4630 3236 4686 3292
rect 4686 3236 4690 3292
rect 4626 3232 4690 3236
rect 11256 3292 11320 3296
rect 11256 3236 11260 3292
rect 11260 3236 11316 3292
rect 11316 3236 11320 3292
rect 11256 3232 11320 3236
rect 11336 3292 11400 3296
rect 11336 3236 11340 3292
rect 11340 3236 11396 3292
rect 11396 3236 11400 3292
rect 11336 3232 11400 3236
rect 11416 3292 11480 3296
rect 11416 3236 11420 3292
rect 11420 3236 11476 3292
rect 11476 3236 11480 3292
rect 11416 3232 11480 3236
rect 11496 3292 11560 3296
rect 11496 3236 11500 3292
rect 11500 3236 11556 3292
rect 11556 3236 11560 3292
rect 11496 3232 11560 3236
rect 18125 3292 18189 3296
rect 18125 3236 18129 3292
rect 18129 3236 18185 3292
rect 18185 3236 18189 3292
rect 18125 3232 18189 3236
rect 18205 3292 18269 3296
rect 18205 3236 18209 3292
rect 18209 3236 18265 3292
rect 18265 3236 18269 3292
rect 18205 3232 18269 3236
rect 18285 3292 18349 3296
rect 18285 3236 18289 3292
rect 18289 3236 18345 3292
rect 18345 3236 18349 3292
rect 18285 3232 18349 3236
rect 18365 3292 18429 3296
rect 18365 3236 18369 3292
rect 18369 3236 18425 3292
rect 18425 3236 18429 3292
rect 18365 3232 18429 3236
rect 7821 2748 7885 2752
rect 7821 2692 7825 2748
rect 7825 2692 7881 2748
rect 7881 2692 7885 2748
rect 7821 2688 7885 2692
rect 7901 2748 7965 2752
rect 7901 2692 7905 2748
rect 7905 2692 7961 2748
rect 7961 2692 7965 2748
rect 7901 2688 7965 2692
rect 7981 2748 8045 2752
rect 7981 2692 7985 2748
rect 7985 2692 8041 2748
rect 8041 2692 8045 2748
rect 7981 2688 8045 2692
rect 8061 2748 8125 2752
rect 8061 2692 8065 2748
rect 8065 2692 8121 2748
rect 8121 2692 8125 2748
rect 8061 2688 8125 2692
rect 14690 2748 14754 2752
rect 14690 2692 14694 2748
rect 14694 2692 14750 2748
rect 14750 2692 14754 2748
rect 14690 2688 14754 2692
rect 14770 2748 14834 2752
rect 14770 2692 14774 2748
rect 14774 2692 14830 2748
rect 14830 2692 14834 2748
rect 14770 2688 14834 2692
rect 14850 2748 14914 2752
rect 14850 2692 14854 2748
rect 14854 2692 14910 2748
rect 14910 2692 14914 2748
rect 14850 2688 14914 2692
rect 14930 2748 14994 2752
rect 14930 2692 14934 2748
rect 14934 2692 14990 2748
rect 14990 2692 14994 2748
rect 14930 2688 14994 2692
rect 4386 2204 4450 2208
rect 4386 2148 4390 2204
rect 4390 2148 4446 2204
rect 4446 2148 4450 2204
rect 4386 2144 4450 2148
rect 4466 2204 4530 2208
rect 4466 2148 4470 2204
rect 4470 2148 4526 2204
rect 4526 2148 4530 2204
rect 4466 2144 4530 2148
rect 4546 2204 4610 2208
rect 4546 2148 4550 2204
rect 4550 2148 4606 2204
rect 4606 2148 4610 2204
rect 4546 2144 4610 2148
rect 4626 2204 4690 2208
rect 4626 2148 4630 2204
rect 4630 2148 4686 2204
rect 4686 2148 4690 2204
rect 4626 2144 4690 2148
rect 11256 2204 11320 2208
rect 11256 2148 11260 2204
rect 11260 2148 11316 2204
rect 11316 2148 11320 2204
rect 11256 2144 11320 2148
rect 11336 2204 11400 2208
rect 11336 2148 11340 2204
rect 11340 2148 11396 2204
rect 11396 2148 11400 2204
rect 11336 2144 11400 2148
rect 11416 2204 11480 2208
rect 11416 2148 11420 2204
rect 11420 2148 11476 2204
rect 11476 2148 11480 2204
rect 11416 2144 11480 2148
rect 11496 2204 11560 2208
rect 11496 2148 11500 2204
rect 11500 2148 11556 2204
rect 11556 2148 11560 2204
rect 11496 2144 11560 2148
rect 18125 2204 18189 2208
rect 18125 2148 18129 2204
rect 18129 2148 18185 2204
rect 18185 2148 18189 2204
rect 18125 2144 18189 2148
rect 18205 2204 18269 2208
rect 18205 2148 18209 2204
rect 18209 2148 18265 2204
rect 18265 2148 18269 2204
rect 18205 2144 18269 2148
rect 18285 2204 18349 2208
rect 18285 2148 18289 2204
rect 18289 2148 18345 2204
rect 18345 2148 18349 2204
rect 18285 2144 18349 2148
rect 18365 2204 18429 2208
rect 18365 2148 18369 2204
rect 18369 2148 18425 2204
rect 18425 2148 18429 2204
rect 18365 2144 18429 2148
<< metal4 >>
rect 4378 21792 4699 22352
rect 4378 21728 4386 21792
rect 4450 21728 4466 21792
rect 4530 21728 4546 21792
rect 4610 21728 4626 21792
rect 4690 21728 4699 21792
rect 4378 20704 4699 21728
rect 4378 20640 4386 20704
rect 4450 20640 4466 20704
rect 4530 20640 4546 20704
rect 4610 20640 4626 20704
rect 4690 20640 4699 20704
rect 4378 19616 4699 20640
rect 4378 19552 4386 19616
rect 4450 19552 4466 19616
rect 4530 19552 4546 19616
rect 4610 19552 4626 19616
rect 4690 19552 4699 19616
rect 4378 19019 4699 19552
rect 4378 18783 4420 19019
rect 4656 18783 4699 19019
rect 4378 18528 4699 18783
rect 4378 18464 4386 18528
rect 4450 18464 4466 18528
rect 4530 18464 4546 18528
rect 4610 18464 4626 18528
rect 4690 18464 4699 18528
rect 4378 17440 4699 18464
rect 4378 17376 4386 17440
rect 4450 17376 4466 17440
rect 4530 17376 4546 17440
rect 4610 17376 4626 17440
rect 4690 17376 4699 17440
rect 4378 16352 4699 17376
rect 4378 16288 4386 16352
rect 4450 16288 4466 16352
rect 4530 16288 4546 16352
rect 4610 16288 4626 16352
rect 4690 16288 4699 16352
rect 4378 15264 4699 16288
rect 4378 15200 4386 15264
rect 4450 15200 4466 15264
rect 4530 15200 4546 15264
rect 4610 15200 4626 15264
rect 4690 15200 4699 15264
rect 4378 14176 4699 15200
rect 4378 14112 4386 14176
rect 4450 14112 4466 14176
rect 4530 14112 4546 14176
rect 4610 14112 4626 14176
rect 4690 14112 4699 14176
rect 4378 13088 4699 14112
rect 4378 13024 4386 13088
rect 4450 13024 4466 13088
rect 4530 13024 4546 13088
rect 4610 13024 4626 13088
rect 4690 13024 4699 13088
rect 4378 12310 4699 13024
rect 4378 12074 4420 12310
rect 4656 12074 4699 12310
rect 4378 12000 4699 12074
rect 4378 11936 4386 12000
rect 4450 11936 4466 12000
rect 4530 11936 4546 12000
rect 4610 11936 4626 12000
rect 4690 11936 4699 12000
rect 4378 10912 4699 11936
rect 4378 10848 4386 10912
rect 4450 10848 4466 10912
rect 4530 10848 4546 10912
rect 4610 10848 4626 10912
rect 4690 10848 4699 10912
rect 4378 9824 4699 10848
rect 4378 9760 4386 9824
rect 4450 9760 4466 9824
rect 4530 9760 4546 9824
rect 4610 9760 4626 9824
rect 4690 9760 4699 9824
rect 4378 8736 4699 9760
rect 4378 8672 4386 8736
rect 4450 8672 4466 8736
rect 4530 8672 4546 8736
rect 4610 8672 4626 8736
rect 4690 8672 4699 8736
rect 4378 7648 4699 8672
rect 4378 7584 4386 7648
rect 4450 7584 4466 7648
rect 4530 7584 4546 7648
rect 4610 7584 4626 7648
rect 4690 7584 4699 7648
rect 4378 6560 4699 7584
rect 4378 6496 4386 6560
rect 4450 6496 4466 6560
rect 4530 6496 4546 6560
rect 4610 6496 4626 6560
rect 4690 6496 4699 6560
rect 4378 5600 4699 6496
rect 4378 5472 4420 5600
rect 4656 5472 4699 5600
rect 4378 5408 4386 5472
rect 4690 5408 4699 5472
rect 4378 5364 4420 5408
rect 4656 5364 4699 5408
rect 4378 4384 4699 5364
rect 4378 4320 4386 4384
rect 4450 4320 4466 4384
rect 4530 4320 4546 4384
rect 4610 4320 4626 4384
rect 4690 4320 4699 4384
rect 4378 3296 4699 4320
rect 4378 3232 4386 3296
rect 4450 3232 4466 3296
rect 4530 3232 4546 3296
rect 4610 3232 4626 3296
rect 4690 3232 4699 3296
rect 4378 2208 4699 3232
rect 4378 2144 4386 2208
rect 4450 2144 4466 2208
rect 4530 2144 4546 2208
rect 4610 2144 4626 2208
rect 4690 2144 4699 2208
rect 4378 2128 4699 2144
rect 7813 22336 8133 22352
rect 7813 22272 7821 22336
rect 7885 22272 7901 22336
rect 7965 22272 7981 22336
rect 8045 22272 8061 22336
rect 8125 22272 8133 22336
rect 7813 21248 8133 22272
rect 7813 21184 7821 21248
rect 7885 21184 7901 21248
rect 7965 21184 7981 21248
rect 8045 21184 8061 21248
rect 8125 21184 8133 21248
rect 7813 20160 8133 21184
rect 7813 20096 7821 20160
rect 7885 20096 7901 20160
rect 7965 20096 7981 20160
rect 8045 20096 8061 20160
rect 8125 20096 8133 20160
rect 7813 19072 8133 20096
rect 7813 19008 7821 19072
rect 7885 19008 7901 19072
rect 7965 19008 7981 19072
rect 8045 19008 8061 19072
rect 8125 19008 8133 19072
rect 7813 17984 8133 19008
rect 7813 17920 7821 17984
rect 7885 17920 7901 17984
rect 7965 17920 7981 17984
rect 8045 17920 8061 17984
rect 8125 17920 8133 17984
rect 7813 16896 8133 17920
rect 7813 16832 7821 16896
rect 7885 16832 7901 16896
rect 7965 16832 7981 16896
rect 8045 16832 8061 16896
rect 8125 16832 8133 16896
rect 7813 15808 8133 16832
rect 7813 15744 7821 15808
rect 7885 15744 7901 15808
rect 7965 15744 7981 15808
rect 8045 15744 8061 15808
rect 8125 15744 8133 15808
rect 7813 15664 8133 15744
rect 7813 15428 7855 15664
rect 8091 15428 8133 15664
rect 7813 14720 8133 15428
rect 7813 14656 7821 14720
rect 7885 14656 7901 14720
rect 7965 14656 7981 14720
rect 8045 14656 8061 14720
rect 8125 14656 8133 14720
rect 7813 13632 8133 14656
rect 7813 13568 7821 13632
rect 7885 13568 7901 13632
rect 7965 13568 7981 13632
rect 8045 13568 8061 13632
rect 8125 13568 8133 13632
rect 7813 12544 8133 13568
rect 7813 12480 7821 12544
rect 7885 12480 7901 12544
rect 7965 12480 7981 12544
rect 8045 12480 8061 12544
rect 8125 12480 8133 12544
rect 7813 11456 8133 12480
rect 7813 11392 7821 11456
rect 7885 11392 7901 11456
rect 7965 11392 7981 11456
rect 8045 11392 8061 11456
rect 8125 11392 8133 11456
rect 7813 10368 8133 11392
rect 7813 10304 7821 10368
rect 7885 10304 7901 10368
rect 7965 10304 7981 10368
rect 8045 10304 8061 10368
rect 8125 10304 8133 10368
rect 7813 9280 8133 10304
rect 7813 9216 7821 9280
rect 7885 9216 7901 9280
rect 7965 9216 7981 9280
rect 8045 9216 8061 9280
rect 8125 9216 8133 9280
rect 7813 8955 8133 9216
rect 7813 8719 7855 8955
rect 8091 8719 8133 8955
rect 7813 8192 8133 8719
rect 7813 8128 7821 8192
rect 7885 8128 7901 8192
rect 7965 8128 7981 8192
rect 8045 8128 8061 8192
rect 8125 8128 8133 8192
rect 7813 7104 8133 8128
rect 7813 7040 7821 7104
rect 7885 7040 7901 7104
rect 7965 7040 7981 7104
rect 8045 7040 8061 7104
rect 8125 7040 8133 7104
rect 7813 6016 8133 7040
rect 7813 5952 7821 6016
rect 7885 5952 7901 6016
rect 7965 5952 7981 6016
rect 8045 5952 8061 6016
rect 8125 5952 8133 6016
rect 7813 4928 8133 5952
rect 7813 4864 7821 4928
rect 7885 4864 7901 4928
rect 7965 4864 7981 4928
rect 8045 4864 8061 4928
rect 8125 4864 8133 4928
rect 7813 3840 8133 4864
rect 7813 3776 7821 3840
rect 7885 3776 7901 3840
rect 7965 3776 7981 3840
rect 8045 3776 8061 3840
rect 8125 3776 8133 3840
rect 7813 2752 8133 3776
rect 7813 2688 7821 2752
rect 7885 2688 7901 2752
rect 7965 2688 7981 2752
rect 8045 2688 8061 2752
rect 8125 2688 8133 2752
rect 7813 2128 8133 2688
rect 11248 21792 11568 22352
rect 11248 21728 11256 21792
rect 11320 21728 11336 21792
rect 11400 21728 11416 21792
rect 11480 21728 11496 21792
rect 11560 21728 11568 21792
rect 11248 20704 11568 21728
rect 11248 20640 11256 20704
rect 11320 20640 11336 20704
rect 11400 20640 11416 20704
rect 11480 20640 11496 20704
rect 11560 20640 11568 20704
rect 11248 19616 11568 20640
rect 11248 19552 11256 19616
rect 11320 19552 11336 19616
rect 11400 19552 11416 19616
rect 11480 19552 11496 19616
rect 11560 19552 11568 19616
rect 11248 19019 11568 19552
rect 11248 18783 11290 19019
rect 11526 18783 11568 19019
rect 11248 18528 11568 18783
rect 11248 18464 11256 18528
rect 11320 18464 11336 18528
rect 11400 18464 11416 18528
rect 11480 18464 11496 18528
rect 11560 18464 11568 18528
rect 11248 17440 11568 18464
rect 11248 17376 11256 17440
rect 11320 17376 11336 17440
rect 11400 17376 11416 17440
rect 11480 17376 11496 17440
rect 11560 17376 11568 17440
rect 11248 16352 11568 17376
rect 11248 16288 11256 16352
rect 11320 16288 11336 16352
rect 11400 16288 11416 16352
rect 11480 16288 11496 16352
rect 11560 16288 11568 16352
rect 11248 15264 11568 16288
rect 11248 15200 11256 15264
rect 11320 15200 11336 15264
rect 11400 15200 11416 15264
rect 11480 15200 11496 15264
rect 11560 15200 11568 15264
rect 11248 14176 11568 15200
rect 11248 14112 11256 14176
rect 11320 14112 11336 14176
rect 11400 14112 11416 14176
rect 11480 14112 11496 14176
rect 11560 14112 11568 14176
rect 11248 13088 11568 14112
rect 11248 13024 11256 13088
rect 11320 13024 11336 13088
rect 11400 13024 11416 13088
rect 11480 13024 11496 13088
rect 11560 13024 11568 13088
rect 11248 12310 11568 13024
rect 11248 12074 11290 12310
rect 11526 12074 11568 12310
rect 11248 12000 11568 12074
rect 11248 11936 11256 12000
rect 11320 11936 11336 12000
rect 11400 11936 11416 12000
rect 11480 11936 11496 12000
rect 11560 11936 11568 12000
rect 11248 10912 11568 11936
rect 11248 10848 11256 10912
rect 11320 10848 11336 10912
rect 11400 10848 11416 10912
rect 11480 10848 11496 10912
rect 11560 10848 11568 10912
rect 11248 9824 11568 10848
rect 11248 9760 11256 9824
rect 11320 9760 11336 9824
rect 11400 9760 11416 9824
rect 11480 9760 11496 9824
rect 11560 9760 11568 9824
rect 11248 8736 11568 9760
rect 11248 8672 11256 8736
rect 11320 8672 11336 8736
rect 11400 8672 11416 8736
rect 11480 8672 11496 8736
rect 11560 8672 11568 8736
rect 11248 7648 11568 8672
rect 11248 7584 11256 7648
rect 11320 7584 11336 7648
rect 11400 7584 11416 7648
rect 11480 7584 11496 7648
rect 11560 7584 11568 7648
rect 11248 6560 11568 7584
rect 11248 6496 11256 6560
rect 11320 6496 11336 6560
rect 11400 6496 11416 6560
rect 11480 6496 11496 6560
rect 11560 6496 11568 6560
rect 11248 5600 11568 6496
rect 11248 5472 11290 5600
rect 11526 5472 11568 5600
rect 11248 5408 11256 5472
rect 11560 5408 11568 5472
rect 11248 5364 11290 5408
rect 11526 5364 11568 5408
rect 11248 4384 11568 5364
rect 11248 4320 11256 4384
rect 11320 4320 11336 4384
rect 11400 4320 11416 4384
rect 11480 4320 11496 4384
rect 11560 4320 11568 4384
rect 11248 3296 11568 4320
rect 11248 3232 11256 3296
rect 11320 3232 11336 3296
rect 11400 3232 11416 3296
rect 11480 3232 11496 3296
rect 11560 3232 11568 3296
rect 11248 2208 11568 3232
rect 11248 2144 11256 2208
rect 11320 2144 11336 2208
rect 11400 2144 11416 2208
rect 11480 2144 11496 2208
rect 11560 2144 11568 2208
rect 11248 2128 11568 2144
rect 14682 22336 15003 22352
rect 14682 22272 14690 22336
rect 14754 22272 14770 22336
rect 14834 22272 14850 22336
rect 14914 22272 14930 22336
rect 14994 22272 15003 22336
rect 14682 21248 15003 22272
rect 14682 21184 14690 21248
rect 14754 21184 14770 21248
rect 14834 21184 14850 21248
rect 14914 21184 14930 21248
rect 14994 21184 15003 21248
rect 14682 20160 15003 21184
rect 14682 20096 14690 20160
rect 14754 20096 14770 20160
rect 14834 20096 14850 20160
rect 14914 20096 14930 20160
rect 14994 20096 15003 20160
rect 14682 19072 15003 20096
rect 14682 19008 14690 19072
rect 14754 19008 14770 19072
rect 14834 19008 14850 19072
rect 14914 19008 14930 19072
rect 14994 19008 15003 19072
rect 14682 17984 15003 19008
rect 14682 17920 14690 17984
rect 14754 17920 14770 17984
rect 14834 17920 14850 17984
rect 14914 17920 14930 17984
rect 14994 17920 15003 17984
rect 14682 16896 15003 17920
rect 14682 16832 14690 16896
rect 14754 16832 14770 16896
rect 14834 16832 14850 16896
rect 14914 16832 14930 16896
rect 14994 16832 15003 16896
rect 14682 15808 15003 16832
rect 14682 15744 14690 15808
rect 14754 15744 14770 15808
rect 14834 15744 14850 15808
rect 14914 15744 14930 15808
rect 14994 15744 15003 15808
rect 14682 15664 15003 15744
rect 14682 15428 14724 15664
rect 14960 15428 15003 15664
rect 14682 14720 15003 15428
rect 14682 14656 14690 14720
rect 14754 14656 14770 14720
rect 14834 14656 14850 14720
rect 14914 14656 14930 14720
rect 14994 14656 15003 14720
rect 14682 13632 15003 14656
rect 14682 13568 14690 13632
rect 14754 13568 14770 13632
rect 14834 13568 14850 13632
rect 14914 13568 14930 13632
rect 14994 13568 15003 13632
rect 14682 12544 15003 13568
rect 14682 12480 14690 12544
rect 14754 12480 14770 12544
rect 14834 12480 14850 12544
rect 14914 12480 14930 12544
rect 14994 12480 15003 12544
rect 14682 11456 15003 12480
rect 14682 11392 14690 11456
rect 14754 11392 14770 11456
rect 14834 11392 14850 11456
rect 14914 11392 14930 11456
rect 14994 11392 15003 11456
rect 14682 10368 15003 11392
rect 14682 10304 14690 10368
rect 14754 10304 14770 10368
rect 14834 10304 14850 10368
rect 14914 10304 14930 10368
rect 14994 10304 15003 10368
rect 14682 9280 15003 10304
rect 14682 9216 14690 9280
rect 14754 9216 14770 9280
rect 14834 9216 14850 9280
rect 14914 9216 14930 9280
rect 14994 9216 15003 9280
rect 14682 8955 15003 9216
rect 14682 8719 14724 8955
rect 14960 8719 15003 8955
rect 14682 8192 15003 8719
rect 14682 8128 14690 8192
rect 14754 8128 14770 8192
rect 14834 8128 14850 8192
rect 14914 8128 14930 8192
rect 14994 8128 15003 8192
rect 14682 7104 15003 8128
rect 14682 7040 14690 7104
rect 14754 7040 14770 7104
rect 14834 7040 14850 7104
rect 14914 7040 14930 7104
rect 14994 7040 15003 7104
rect 14682 6016 15003 7040
rect 14682 5952 14690 6016
rect 14754 5952 14770 6016
rect 14834 5952 14850 6016
rect 14914 5952 14930 6016
rect 14994 5952 15003 6016
rect 14682 4928 15003 5952
rect 14682 4864 14690 4928
rect 14754 4864 14770 4928
rect 14834 4864 14850 4928
rect 14914 4864 14930 4928
rect 14994 4864 15003 4928
rect 14682 3840 15003 4864
rect 14682 3776 14690 3840
rect 14754 3776 14770 3840
rect 14834 3776 14850 3840
rect 14914 3776 14930 3840
rect 14994 3776 15003 3840
rect 14682 2752 15003 3776
rect 14682 2688 14690 2752
rect 14754 2688 14770 2752
rect 14834 2688 14850 2752
rect 14914 2688 14930 2752
rect 14994 2688 15003 2752
rect 14682 2128 15003 2688
rect 18117 21792 18437 22352
rect 18117 21728 18125 21792
rect 18189 21728 18205 21792
rect 18269 21728 18285 21792
rect 18349 21728 18365 21792
rect 18429 21728 18437 21792
rect 18117 20704 18437 21728
rect 18117 20640 18125 20704
rect 18189 20640 18205 20704
rect 18269 20640 18285 20704
rect 18349 20640 18365 20704
rect 18429 20640 18437 20704
rect 18117 19616 18437 20640
rect 18117 19552 18125 19616
rect 18189 19552 18205 19616
rect 18269 19552 18285 19616
rect 18349 19552 18365 19616
rect 18429 19552 18437 19616
rect 18117 19019 18437 19552
rect 18117 18783 18159 19019
rect 18395 18783 18437 19019
rect 18117 18528 18437 18783
rect 18117 18464 18125 18528
rect 18189 18464 18205 18528
rect 18269 18464 18285 18528
rect 18349 18464 18365 18528
rect 18429 18464 18437 18528
rect 18117 17440 18437 18464
rect 18117 17376 18125 17440
rect 18189 17376 18205 17440
rect 18269 17376 18285 17440
rect 18349 17376 18365 17440
rect 18429 17376 18437 17440
rect 18117 16352 18437 17376
rect 18117 16288 18125 16352
rect 18189 16288 18205 16352
rect 18269 16288 18285 16352
rect 18349 16288 18365 16352
rect 18429 16288 18437 16352
rect 18117 15264 18437 16288
rect 18117 15200 18125 15264
rect 18189 15200 18205 15264
rect 18269 15200 18285 15264
rect 18349 15200 18365 15264
rect 18429 15200 18437 15264
rect 18117 14176 18437 15200
rect 18117 14112 18125 14176
rect 18189 14112 18205 14176
rect 18269 14112 18285 14176
rect 18349 14112 18365 14176
rect 18429 14112 18437 14176
rect 18117 13088 18437 14112
rect 18117 13024 18125 13088
rect 18189 13024 18205 13088
rect 18269 13024 18285 13088
rect 18349 13024 18365 13088
rect 18429 13024 18437 13088
rect 18117 12310 18437 13024
rect 18117 12074 18159 12310
rect 18395 12074 18437 12310
rect 18117 12000 18437 12074
rect 18117 11936 18125 12000
rect 18189 11936 18205 12000
rect 18269 11936 18285 12000
rect 18349 11936 18365 12000
rect 18429 11936 18437 12000
rect 18117 10912 18437 11936
rect 18117 10848 18125 10912
rect 18189 10848 18205 10912
rect 18269 10848 18285 10912
rect 18349 10848 18365 10912
rect 18429 10848 18437 10912
rect 18117 9824 18437 10848
rect 18117 9760 18125 9824
rect 18189 9760 18205 9824
rect 18269 9760 18285 9824
rect 18349 9760 18365 9824
rect 18429 9760 18437 9824
rect 18117 8736 18437 9760
rect 18117 8672 18125 8736
rect 18189 8672 18205 8736
rect 18269 8672 18285 8736
rect 18349 8672 18365 8736
rect 18429 8672 18437 8736
rect 18117 7648 18437 8672
rect 18117 7584 18125 7648
rect 18189 7584 18205 7648
rect 18269 7584 18285 7648
rect 18349 7584 18365 7648
rect 18429 7584 18437 7648
rect 18117 6560 18437 7584
rect 18117 6496 18125 6560
rect 18189 6496 18205 6560
rect 18269 6496 18285 6560
rect 18349 6496 18365 6560
rect 18429 6496 18437 6560
rect 18117 5600 18437 6496
rect 18117 5472 18159 5600
rect 18395 5472 18437 5600
rect 18117 5408 18125 5472
rect 18429 5408 18437 5472
rect 18117 5364 18159 5408
rect 18395 5364 18437 5408
rect 18117 4384 18437 5364
rect 18117 4320 18125 4384
rect 18189 4320 18205 4384
rect 18269 4320 18285 4384
rect 18349 4320 18365 4384
rect 18429 4320 18437 4384
rect 18117 3296 18437 4320
rect 18117 3232 18125 3296
rect 18189 3232 18205 3296
rect 18269 3232 18285 3296
rect 18349 3232 18365 3296
rect 18429 3232 18437 3296
rect 18117 2208 18437 3232
rect 18117 2144 18125 2208
rect 18189 2144 18205 2208
rect 18269 2144 18285 2208
rect 18349 2144 18365 2208
rect 18429 2144 18437 2208
rect 18117 2128 18437 2144
<< via4 >>
rect 4420 18783 4656 19019
rect 4420 12074 4656 12310
rect 4420 5472 4656 5600
rect 4420 5408 4450 5472
rect 4450 5408 4466 5472
rect 4466 5408 4530 5472
rect 4530 5408 4546 5472
rect 4546 5408 4610 5472
rect 4610 5408 4626 5472
rect 4626 5408 4656 5472
rect 4420 5364 4656 5408
rect 7855 15428 8091 15664
rect 7855 8719 8091 8955
rect 11290 18783 11526 19019
rect 11290 12074 11526 12310
rect 11290 5472 11526 5600
rect 11290 5408 11320 5472
rect 11320 5408 11336 5472
rect 11336 5408 11400 5472
rect 11400 5408 11416 5472
rect 11416 5408 11480 5472
rect 11480 5408 11496 5472
rect 11496 5408 11526 5472
rect 11290 5364 11526 5408
rect 14724 15428 14960 15664
rect 14724 8719 14960 8955
rect 18159 18783 18395 19019
rect 18159 12074 18395 12310
rect 18159 5472 18395 5600
rect 18159 5408 18189 5472
rect 18189 5408 18205 5472
rect 18205 5408 18269 5472
rect 18269 5408 18285 5472
rect 18285 5408 18349 5472
rect 18349 5408 18365 5472
rect 18365 5408 18395 5472
rect 18159 5364 18395 5408
<< metal5 >>
rect 1104 19019 21712 19061
rect 1104 18783 4420 19019
rect 4656 18783 11290 19019
rect 11526 18783 18159 19019
rect 18395 18783 21712 19019
rect 1104 18741 21712 18783
rect 1104 15664 21712 15707
rect 1104 15428 7855 15664
rect 8091 15428 14724 15664
rect 14960 15428 21712 15664
rect 1104 15386 21712 15428
rect 1104 12310 21712 12352
rect 1104 12074 4420 12310
rect 4656 12074 11290 12310
rect 11526 12074 18159 12310
rect 18395 12074 21712 12310
rect 1104 12032 21712 12074
rect 1104 8955 21712 8997
rect 1104 8719 7855 8955
rect 8091 8719 14724 8955
rect 14960 8719 21712 8955
rect 1104 8677 21712 8719
rect 1104 5600 21712 5643
rect 1104 5364 4420 5600
rect 4656 5364 11290 5600
rect 11526 5364 18159 5600
rect 18395 5364 21712 5600
rect 1104 5322 21712 5364
use sky130_fd_sc_hd__decap_8  FILLER_1_16
timestamp 1616762085
transform 1 0 2576 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_11
timestamp 1616762085
transform 1 0 2116 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1616762085
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_12
timestamp 1616762085
transform 1 0 2208 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3
timestamp 1616762085
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_38
timestamp 1616762085
transform 1 0 2208 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1616762085
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1616762085
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _51_
timestamp 1616762085
transform 1 0 1932 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1616762085
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1616762085
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30
timestamp 1616762085
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24
timestamp 1616762085
transform 1 0 3312 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1616762085
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _52_
timestamp 1616762085
transform 1 0 3312 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1616762085
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1616762085
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1616762085
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1616762085
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51
timestamp 1616762085
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1616762085
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1616762085
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1616762085
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1616762085
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1616762085
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1616762085
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1616762085
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1616762085
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1616762085
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1616762085
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1616762085
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1616762085
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1616762085
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1616762085
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1616762085
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1616762085
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1616762085
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1616762085
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1616762085
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1616762085
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1616762085
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1616762085
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1616762085
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1616762085
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1616762085
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1616762085
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1616762085
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1616762085
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1616762085
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1616762085
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1616762085
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1616762085
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1616762085
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1616762085
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1616762085
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_218
timestamp 1616762085
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1616762085
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1616762085
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_220
timestamp 1616762085
transform 1 0 21344 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1616762085
transform -1 0 21712 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1616762085
transform -1 0 21712 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_16
timestamp 1616762085
transform 1 0 2576 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_11
timestamp 1616762085
transform 1 0 2116 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1616762085
transform 1 0 1380 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_28
timestamp 1616762085
transform 1 0 2208 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1616762085
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_32
timestamp 1616762085
transform 1 0 4048 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1616762085
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1616762085
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1616762085
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_34
timestamp 1616762085
transform 1 0 4784 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1616762085
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1616762085
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1616762085
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1616762085
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1616762085
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1616762085
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1616762085
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1616762085
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1616762085
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1616762085
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1616762085
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1616762085
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1616762085
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1616762085
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1616762085
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_215
timestamp 1616762085
transform 1 0 20884 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1616762085
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1616762085
transform -1 0 21712 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_16
timestamp 1616762085
transform 1 0 2576 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1616762085
transform 1 0 2116 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1616762085
transform 1 0 1380 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_18
timestamp 1616762085
transform 1 0 2208 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1616762085
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_28
timestamp 1616762085
transform 1 0 3680 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_35
timestamp 1616762085
transform 1 0 3312 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1616762085
transform 1 0 5152 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_17
timestamp 1616762085
transform 1 0 4784 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1616762085
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1616762085
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_56
timestamp 1616762085
transform 1 0 6256 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1616762085
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1616762085
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1616762085
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1616762085
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1616762085
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1616762085
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1616762085
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1616762085
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1616762085
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1616762085
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1616762085
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1616762085
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1616762085
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1616762085
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1616762085
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_220
timestamp 1616762085
transform 1 0 21344 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1616762085
transform -1 0 21712 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_16
timestamp 1616762085
transform 1 0 2576 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1616762085
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1616762085
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _53_
timestamp 1616762085
transform 1 0 1472 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1616762085
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1616762085
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1616762085
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_43
timestamp 1616762085
transform 1 0 5060 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _27_
timestamp 1616762085
transform 1 0 4416 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_4_67
timestamp 1616762085
transform 1 0 7268 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_55
timestamp 1616762085
transform 1 0 6164 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_36
timestamp 1616762085
transform 1 0 6900 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_22
timestamp 1616762085
transform 1 0 5796 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_79
timestamp 1616762085
transform 1 0 8372 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1616762085
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1616762085
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1616762085
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1616762085
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1616762085
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1616762085
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1616762085
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1616762085
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1616762085
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1616762085
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1616762085
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1616762085
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1616762085
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_215
timestamp 1616762085
transform 1 0 20884 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1616762085
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1616762085
transform -1 0 21712 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1616762085
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1616762085
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _54_
timestamp 1616762085
transform 1 0 1932 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_25
timestamp 1616762085
transform 1 0 3404 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _55_
timestamp 1616762085
transform 1 0 4140 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_5_49
timestamp 1616762085
transform 1 0 5612 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_66
timestamp 1616762085
transform 1 0 7176 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_27
timestamp 1616762085
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1616762085
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_78
timestamp 1616762085
transform 1 0 8280 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_90
timestamp 1616762085
transform 1 0 9384 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_114
timestamp 1616762085
transform 1 0 11592 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_102
timestamp 1616762085
transform 1 0 10488 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1616762085
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1616762085
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1616762085
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1616762085
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1616762085
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1616762085
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1616762085
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1616762085
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1616762085
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1616762085
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_220
timestamp 1616762085
transform 1 0 21344 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1616762085
transform -1 0 21712 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_14
timestamp 1616762085
transform 1 0 2392 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1616762085
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1616762085
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1616762085
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _29_
timestamp 1616762085
transform 1 0 1380 0 -1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _28_
timestamp 1616762085
transform 1 0 1748 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_7_26
timestamp 1616762085
transform 1 0 3496 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_32
timestamp 1616762085
transform 1 0 4048 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1616762085
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_17
timestamp 1616762085
transform 1 0 2668 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1616762085
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _30_
timestamp 1616762085
transform 1 0 4048 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_7_46
timestamp 1616762085
transform 1 0 5336 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _56_
timestamp 1616762085
transform 1 0 4784 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1616762085
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1616762085
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1616762085
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1616762085
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _31_
timestamp 1616762085
transform 1 0 6900 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_7_77
timestamp 1616762085
transform 1 0 8188 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_75
timestamp 1616762085
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_68
timestamp 1616762085
transform 1 0 7360 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_4
timestamp 1616762085
transform 1 0 7636 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_101
timestamp 1616762085
transform 1 0 10396 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_89
timestamp 1616762085
transform 1 0 9292 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1616762085
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1616762085
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1616762085
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1616762085
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1616762085
transform 1 0 11500 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1616762085
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1616762085
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1616762085
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1616762085
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1616762085
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1616762085
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1616762085
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1616762085
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1616762085
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1616762085
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1616762085
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1616762085
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1616762085
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1616762085
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1616762085
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1616762085
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1616762085
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1616762085
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1616762085
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1616762085
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1616762085
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_215
timestamp 1616762085
transform 1 0 20884 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1616762085
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_220
timestamp 1616762085
transform 1 0 21344 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1616762085
transform -1 0 21712 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1616762085
transform -1 0 21712 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_16
timestamp 1616762085
transform 1 0 2576 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_11
timestamp 1616762085
transform 1 0 2116 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1616762085
transform 1 0 1380 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_6
timestamp 1616762085
transform 1 0 2208 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1616762085
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_32
timestamp 1616762085
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_28
timestamp 1616762085
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1616762085
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_44
timestamp 1616762085
transform 1 0 5152 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_5
timestamp 1616762085
transform 1 0 4784 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_56
timestamp 1616762085
transform 1 0 6256 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_10
timestamp 1616762085
transform 1 0 5888 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _57_
timestamp 1616762085
transform 1 0 6992 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1616762085
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1616762085
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1616762085
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1616762085
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1616762085
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1616762085
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1616762085
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1616762085
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1616762085
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1616762085
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1616762085
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1616762085
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1616762085
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_215
timestamp 1616762085
transform 1 0 20884 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1616762085
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1616762085
transform -1 0 21712 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_16
timestamp 1616762085
transform 1 0 2576 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_11
timestamp 1616762085
transform 1 0 2116 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1616762085
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_12
timestamp 1616762085
transform 1 0 2208 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1616762085
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_28
timestamp 1616762085
transform 1 0 3680 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_32
timestamp 1616762085
transform 1 0 3312 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_44
timestamp 1616762085
transform 1 0 5152 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_11
timestamp 1616762085
transform 1 0 4784 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1616762085
transform 1 0 6808 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1616762085
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_56
timestamp 1616762085
transform 1 0 6256 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1616762085
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_70
timestamp 1616762085
transform 1 0 7544 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _58_
timestamp 1616762085
transform 1 0 7636 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_99
timestamp 1616762085
transform 1 0 10212 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_87
timestamp 1616762085
transform 1 0 9108 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_21
timestamp 1616762085
transform 1 0 9844 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_111
timestamp 1616762085
transform 1 0 11316 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1616762085
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp 1616762085
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1616762085
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1616762085
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1616762085
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1616762085
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1616762085
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1616762085
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1616762085
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1616762085
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1616762085
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_220
timestamp 1616762085
transform 1 0 21344 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1616762085
transform -1 0 21712 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_16
timestamp 1616762085
transform 1 0 2576 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1616762085
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1616762085
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_23
timestamp 1616762085
transform 1 0 2208 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1616762085
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_32
timestamp 1616762085
transform 1 0 4048 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_28
timestamp 1616762085
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1616762085
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_44
timestamp 1616762085
transform 1 0 5152 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_31
timestamp 1616762085
transform 1 0 4784 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_59
timestamp 1616762085
transform 1 0 6532 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_52
timestamp 1616762085
transform 1 0 5888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_30
timestamp 1616762085
transform 1 0 6164 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _26_
timestamp 1616762085
transform 1 0 7268 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_10_74
timestamp 1616762085
transform 1 0 7912 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1616762085
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_86
timestamp 1616762085
transform 1 0 9016 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1616762085
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1616762085
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1616762085
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1616762085
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1616762085
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1616762085
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1616762085
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1616762085
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1616762085
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1616762085
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1616762085
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_215
timestamp 1616762085
transform 1 0 20884 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1616762085
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1616762085
transform -1 0 21712 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_16
timestamp 1616762085
transform 1 0 2576 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_11
timestamp 1616762085
transform 1 0 2116 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1616762085
transform 1 0 1380 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_37
timestamp 1616762085
transform 1 0 2208 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1616762085
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_28
timestamp 1616762085
transform 1 0 3680 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_40
timestamp 1616762085
transform 1 0 4784 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_62
timestamp 1616762085
transform 1 0 6808 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1616762085
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_52
timestamp 1616762085
transform 1 0 5888 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1616762085
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_75
timestamp 1616762085
transform 1 0 8004 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_70
timestamp 1616762085
transform 1 0 7544 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_33
timestamp 1616762085
transform 1 0 8740 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_16
timestamp 1616762085
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_99
timestamp 1616762085
transform 1 0 10212 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_87
timestamp 1616762085
transform 1 0 9108 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_106
timestamp 1616762085
transform 1 0 10856 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_3
timestamp 1616762085
transform 1 0 10488 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1616762085
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1616762085
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1616762085
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1616762085
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1616762085
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1616762085
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1616762085
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1616762085
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1616762085
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1616762085
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1616762085
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_220
timestamp 1616762085
transform 1 0 21344 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1616762085
transform -1 0 21712 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1616762085
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1616762085
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1616762085
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1616762085
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1616762085
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1616762085
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1616762085
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1616762085
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_75
timestamp 1616762085
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_68
timestamp 1616762085
transform 1 0 7360 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_26
timestamp 1616762085
transform 1 0 7636 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1616762085
transform 1 0 9660 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1616762085
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1616762085
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1616762085
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _35_
timestamp 1616762085
transform 1 0 9752 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_12_108
timestamp 1616762085
transform 1 0 11040 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_132
timestamp 1616762085
transform 1 0 13248 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_120
timestamp 1616762085
transform 1 0 12144 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_144
timestamp 1616762085
transform 1 0 14352 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1616762085
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1616762085
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1616762085
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1616762085
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1616762085
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1616762085
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1616762085
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_215
timestamp 1616762085
transform 1 0 20884 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1616762085
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1616762085
transform -1 0 21712 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1616762085
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1616762085
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1616762085
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1616762085
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1616762085
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1616762085
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1616762085
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1616762085
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1616762085
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1616762085
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1616762085
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1616762085
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1616762085
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1616762085
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1616762085
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1616762085
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1616762085
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1616762085
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1616762085
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1616762085
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_101
timestamp 1616762085
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_93
timestamp 1616762085
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_94
timestamp 1616762085
transform 1 0 9752 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_86
timestamp 1616762085
transform 1 0 9016 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1616762085
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _25_
timestamp 1616762085
transform 1 0 9844 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_13_111
timestamp 1616762085
transform 1 0 11316 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _32_
timestamp 1616762085
transform 1 0 10580 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_131
timestamp 1616762085
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_119
timestamp 1616762085
transform 1 0 12052 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1616762085
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1616762085
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_15
timestamp 1616762085
transform 1 0 12788 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1616762085
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1616762085
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_143
timestamp 1616762085
transform 1 0 14260 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1616762085
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1616762085
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1616762085
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1616762085
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1616762085
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1616762085
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1616762085
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1616762085
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1616762085
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1616762085
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1616762085
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1616762085
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1616762085
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_215
timestamp 1616762085
transform 1 0 20884 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1616762085
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1616762085
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_220
timestamp 1616762085
transform 1 0 21344 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1616762085
transform -1 0 21712 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1616762085
transform -1 0 21712 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1616762085
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1616762085
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1616762085
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1616762085
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1616762085
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1616762085
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1616762085
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1616762085
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1616762085
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1616762085
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_90
timestamp 1616762085
transform 1 0 9384 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_25
timestamp 1616762085
transform 1 0 9016 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _34_
timestamp 1616762085
transform 1 0 10120 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_15_117
timestamp 1616762085
transform 1 0 11868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_105
timestamp 1616762085
transform 1 0 10764 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1616762085
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1616762085
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1616762085
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1616762085
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1616762085
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_159
timestamp 1616762085
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1616762085
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_171
timestamp 1616762085
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1616762085
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1616762085
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1616762085
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_220
timestamp 1616762085
transform 1 0 21344 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1616762085
transform -1 0 21712 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1616762085
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1616762085
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1616762085
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1616762085
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1616762085
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1616762085
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1616762085
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1616762085
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1616762085
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1616762085
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 1616762085
transform 1 0 10396 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1616762085
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1616762085
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_106
timestamp 1616762085
transform 1 0 10856 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_29
timestamp 1616762085
transform 1 0 11592 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_9
timestamp 1616762085
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_130
timestamp 1616762085
transform 1 0 13064 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_118
timestamp 1616762085
transform 1 0 11960 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_24
timestamp 1616762085
transform 1 0 13340 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1616762085
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_137
timestamp 1616762085
transform 1 0 13708 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1616762085
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1616762085
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1616762085
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1616762085
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1616762085
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1616762085
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_215
timestamp 1616762085
transform 1 0 20884 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1616762085
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1616762085
transform -1 0 21712 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1616762085
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1616762085
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1616762085
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1616762085
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1616762085
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1616762085
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1616762085
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1616762085
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1616762085
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1616762085
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_98
timestamp 1616762085
transform 1 0 10120 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1616762085
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_106
timestamp 1616762085
transform 1 0 10856 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_20
timestamp 1616762085
transform 1 0 10488 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1616762085
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_123
timestamp 1616762085
transform 1 0 12420 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1616762085
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_2
timestamp 1616762085
transform 1 0 13340 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1616762085
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1616762085
transform 1 0 14812 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1616762085
transform 1 0 13708 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_161
timestamp 1616762085
transform 1 0 15916 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1616762085
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1616762085
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_173
timestamp 1616762085
transform 1 0 17020 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1616762085
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1616762085
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1616762085
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_220
timestamp 1616762085
transform 1 0 21344 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1616762085
transform -1 0 21712 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1616762085
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1616762085
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1616762085
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1616762085
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1616762085
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1616762085
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1616762085
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1616762085
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1616762085
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1616762085
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1616762085
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1616762085
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_117
timestamp 1616762085
transform 1 0 11868 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1616762085
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_125
timestamp 1616762085
transform 1 0 12604 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _33_
timestamp 1616762085
transform 1 0 12696 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1616762085
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_142
timestamp 1616762085
transform 1 0 14168 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1616762085
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1616762085
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1616762085
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1616762085
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1616762085
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1616762085
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_215
timestamp 1616762085
transform 1 0 20884 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1616762085
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1616762085
transform -1 0 21712 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1616762085
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1616762085
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1616762085
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1616762085
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1616762085
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1616762085
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1616762085
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1616762085
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1616762085
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1616762085
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1616762085
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1616762085
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1616762085
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1616762085
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1616762085
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1616762085
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1616762085
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1616762085
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1616762085
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1616762085
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1616762085
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1616762085
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1616762085
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1616762085
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_117
timestamp 1616762085
transform 1 0 11868 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1616762085
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1616762085
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_131
timestamp 1616762085
transform 1 0 13156 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_123
timestamp 1616762085
transform 1 0 12420 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1616762085
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _39_
timestamp 1616762085
transform 1 0 12604 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__a2bb2o_4  _36_
timestamp 1616762085
transform 1 0 13432 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1616762085
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_139
timestamp 1616762085
transform 1 0 13892 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_150
timestamp 1616762085
transform 1 0 14904 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1616762085
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1616762085
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_162
timestamp 1616762085
transform 1 0 16008 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_8
timestamp 1616762085
transform 1 0 15640 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1616762085
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1616762085
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1616762085
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1616762085
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_174
timestamp 1616762085
transform 1 0 17112 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1616762085
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1616762085
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1616762085
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1616762085
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_215
timestamp 1616762085
transform 1 0 20884 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1616762085
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1616762085
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_220
timestamp 1616762085
transform 1 0 21344 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1616762085
transform -1 0 21712 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1616762085
transform -1 0 21712 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1616762085
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1616762085
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1616762085
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1616762085
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1616762085
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1616762085
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1616762085
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1616762085
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1616762085
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1616762085
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1616762085
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1616762085
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1616762085
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_123
timestamp 1616762085
transform 1 0 12420 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1616762085
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _38_
timestamp 1616762085
transform 1 0 12972 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_21_148
timestamp 1616762085
transform 1 0 14720 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_136
timestamp 1616762085
transform 1 0 13616 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_19
timestamp 1616762085
transform 1 0 14352 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_160
timestamp 1616762085
transform 1 0 15824 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1616762085
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_180
timestamp 1616762085
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_172
timestamp 1616762085
transform 1 0 16928 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1616762085
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1616762085
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1616762085
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_220
timestamp 1616762085
transform 1 0 21344 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1616762085
transform -1 0 21712 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1616762085
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1616762085
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1616762085
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1616762085
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1616762085
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1616762085
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1616762085
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1616762085
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1616762085
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1616762085
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1616762085
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1616762085
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1616762085
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1616762085
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_129
timestamp 1616762085
transform 1 0 12972 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_14
timestamp 1616762085
transform 1 0 13340 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1616762085
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1616762085
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_162
timestamp 1616762085
transform 1 0 16008 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_154
timestamp 1616762085
transform 1 0 15272 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1616762085
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _40_
timestamp 1616762085
transform 1 0 16284 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_22_181
timestamp 1616762085
transform 1 0 17756 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_193
timestamp 1616762085
transform 1 0 18860 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_215
timestamp 1616762085
transform 1 0 20884 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_213
timestamp 1616762085
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_205
timestamp 1616762085
transform 1 0 19964 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1616762085
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1616762085
transform -1 0 21712 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1616762085
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1616762085
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1616762085
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1616762085
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1616762085
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1616762085
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1616762085
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1616762085
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1616762085
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1616762085
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1616762085
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1616762085
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1616762085
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1616762085
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1616762085
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1616762085
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1616762085
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_167
timestamp 1616762085
transform 1 0 16468 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_159
timestamp 1616762085
transform 1 0 15732 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _42_
timestamp 1616762085
transform 1 0 15824 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1616762085
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1616762085
transform 1 0 17572 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1616762085
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1616762085
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1616762085
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_220
timestamp 1616762085
transform 1 0 21344 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1616762085
transform -1 0 21712 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1616762085
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1616762085
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1616762085
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1616762085
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1616762085
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1616762085
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1616762085
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1616762085
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1616762085
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1616762085
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1616762085
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1616762085
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1616762085
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1616762085
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1616762085
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1616762085
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1616762085
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1616762085
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _37_
timestamp 1616762085
transform 1 0 15548 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_185
timestamp 1616762085
transform 1 0 18124 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_173
timestamp 1616762085
transform 1 0 17020 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_1
timestamp 1616762085
transform 1 0 17756 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1616762085
transform 1 0 19228 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_13
timestamp 1616762085
transform 1 0 18860 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_215
timestamp 1616762085
transform 1 0 20884 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1616762085
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1616762085
transform 1 0 20332 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1616762085
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1616762085
transform -1 0 21712 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1616762085
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1616762085
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1616762085
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1616762085
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1616762085
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1616762085
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1616762085
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1616762085
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1616762085
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1616762085
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1616762085
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1616762085
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1616762085
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1616762085
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1616762085
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_147
timestamp 1616762085
transform 1 0 14628 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1616762085
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_155
timestamp 1616762085
transform 1 0 15364 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _43_
timestamp 1616762085
transform 1 0 15456 0 1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1616762085
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1616762085
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_170
timestamp 1616762085
transform 1 0 16744 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1616762085
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1616762085
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1616762085
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_220
timestamp 1616762085
transform 1 0 21344 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1616762085
transform -1 0 21712 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1616762085
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1616762085
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1616762085
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1616762085
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1616762085
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1616762085
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1616762085
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1616762085
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1616762085
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1616762085
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1616762085
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1616762085
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1616762085
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1616762085
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1616762085
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1616762085
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1616762085
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1616762085
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1616762085
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1616762085
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1616762085
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1616762085
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1616762085
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1616762085
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1616762085
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1616762085
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1616762085
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1616762085
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1616762085
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1616762085
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1616762085
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1616762085
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1616762085
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1616762085
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1616762085
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_162
timestamp 1616762085
transform 1 0 16008 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_154
timestamp 1616762085
transform 1 0 15272 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_7
timestamp 1616762085
transform 1 0 16192 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1616762085
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1616762085
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1616762085
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_180
timestamp 1616762085
transform 1 0 17664 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1616762085
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_201
timestamp 1616762085
transform 1 0 19596 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_196
timestamp 1616762085
transform 1 0 19136 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_192
timestamp 1616762085
transform 1 0 18768 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_0
timestamp 1616762085
transform 1 0 19228 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_213
timestamp 1616762085
transform 1 0 20700 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_215
timestamp 1616762085
transform 1 0 20884 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1616762085
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_204
timestamp 1616762085
transform 1 0 19872 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1616762085
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1616762085
transform -1 0 21712 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1616762085
transform -1 0 21712 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1616762085
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1616762085
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1616762085
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1616762085
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1616762085
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1616762085
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1616762085
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1616762085
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1616762085
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1616762085
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1616762085
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1616762085
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1616762085
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1616762085
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1616762085
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1616762085
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1616762085
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1616762085
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1616762085
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1616762085
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _44_
timestamp 1616762085
transform 1 0 18584 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_28_215
timestamp 1616762085
transform 1 0 20884 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_206
timestamp 1616762085
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1616762085
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1616762085
transform -1 0 21712 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1616762085
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1616762085
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1616762085
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1616762085
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1616762085
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1616762085
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1616762085
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1616762085
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1616762085
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1616762085
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1616762085
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1616762085
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1616762085
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1616762085
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1616762085
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1616762085
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1616762085
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1616762085
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_184
timestamp 1616762085
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1616762085
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1616762085
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _41_
timestamp 1616762085
transform 1 0 18584 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_29_218
timestamp 1616762085
transform 1 0 21160 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_206
timestamp 1616762085
transform 1 0 20056 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1616762085
transform -1 0 21712 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1616762085
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1616762085
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1616762085
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1616762085
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1616762085
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1616762085
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1616762085
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1616762085
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1616762085
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1616762085
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1616762085
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1616762085
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1616762085
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1616762085
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1616762085
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1616762085
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1616762085
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1616762085
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1616762085
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1616762085
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _47_
timestamp 1616762085
transform 1 0 18584 0 -1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_30_215
timestamp 1616762085
transform 1 0 20884 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1616762085
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_204
timestamp 1616762085
transform 1 0 19872 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1616762085
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1616762085
transform -1 0 21712 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1616762085
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1616762085
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1616762085
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1616762085
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1616762085
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1616762085
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1616762085
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1616762085
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1616762085
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1616762085
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1616762085
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1616762085
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1616762085
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1616762085
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1616762085
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1616762085
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1616762085
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1616762085
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_184
timestamp 1616762085
transform 1 0 18032 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1616762085
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1616762085
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_200
timestamp 1616762085
transform 1 0 19504 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_192
timestamp 1616762085
transform 1 0 18768 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _46_
timestamp 1616762085
transform 1 0 18860 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_31_212
timestamp 1616762085
transform 1 0 20608 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_220
timestamp 1616762085
transform 1 0 21344 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1616762085
transform -1 0 21712 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1616762085
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1616762085
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1616762085
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1616762085
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1616762085
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1616762085
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1616762085
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1616762085
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1616762085
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1616762085
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1616762085
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1616762085
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1616762085
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1616762085
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1616762085
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1616762085
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1616762085
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1616762085
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1616762085
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1616762085
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_198
timestamp 1616762085
transform 1 0 19320 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_190
timestamp 1616762085
transform 1 0 18584 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _45_
timestamp 1616762085
transform 1 0 19412 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_32_215
timestamp 1616762085
transform 1 0 20884 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_206
timestamp 1616762085
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1616762085
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1616762085
transform -1 0 21712 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1616762085
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1616762085
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1616762085
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1616762085
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1616762085
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1616762085
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1616762085
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1616762085
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1616762085
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1616762085
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1616762085
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1616762085
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1616762085
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1616762085
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1616762085
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1616762085
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1616762085
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1616762085
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1616762085
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1616762085
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1616762085
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1616762085
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1616762085
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1616762085
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1616762085
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1616762085
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1616762085
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1616762085
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1616762085
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1616762085
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1616762085
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1616762085
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1616762085
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1616762085
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1616762085
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1616762085
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1616762085
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1616762085
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1616762085
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1616762085
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1616762085
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_190
timestamp 1616762085
transform 1 0 18584 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_196
timestamp 1616762085
transform 1 0 19136 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _49_
timestamp 1616762085
transform 1 0 19228 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _48_
timestamp 1616762085
transform 1 0 18768 0 -1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_34_215
timestamp 1616762085
transform 1 0 20884 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_206
timestamp 1616762085
transform 1 0 20056 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_213
timestamp 1616762085
transform 1 0 20700 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1616762085
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1616762085
transform -1 0 21712 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1616762085
transform -1 0 21712 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1616762085
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1616762085
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1616762085
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1616762085
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1616762085
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1616762085
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1616762085
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1616762085
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1616762085
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1616762085
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1616762085
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1616762085
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_110
timestamp 1616762085
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1616762085
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1616762085
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1616762085
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1616762085
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1616762085
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1616762085
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1616762085
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1616762085
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_196
timestamp 1616762085
transform 1 0 19136 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _50_
timestamp 1616762085
transform 1 0 19228 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_35_213
timestamp 1616762085
transform 1 0 20700 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1616762085
transform -1 0 21712 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1616762085
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1616762085
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1616762085
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1616762085
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1616762085
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1616762085
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1616762085
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_63
timestamp 1616762085
transform 1 0 6900 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_56
timestamp 1616762085
transform 1 0 6256 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1616762085
transform 1 0 6808 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_75
timestamp 1616762085
transform 1 0 8004 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_94
timestamp 1616762085
transform 1 0 9752 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_87
timestamp 1616762085
transform 1 0 9108 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1616762085
transform 1 0 9660 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_106
timestamp 1616762085
transform 1 0 10856 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_125
timestamp 1616762085
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_118
timestamp 1616762085
transform 1 0 11960 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1616762085
transform 1 0 12512 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_149
timestamp 1616762085
transform 1 0 14812 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_137
timestamp 1616762085
transform 1 0 13708 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1616762085
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1616762085
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1616762085
transform 1 0 15364 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_180
timestamp 1616762085
transform 1 0 17664 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_199
timestamp 1616762085
transform 1 0 19412 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_187
timestamp 1616762085
transform 1 0 18308 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1616762085
transform 1 0 18216 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_218
timestamp 1616762085
transform 1 0 21160 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_211
timestamp 1616762085
transform 1 0 20516 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1616762085
transform 1 0 21068 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1616762085
transform -1 0 21712 0 -1 22304
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 12520 800 12640 4 ci
port 1 nsew
rlabel metal3 s 22058 23536 22858 23656 4 co
port 2 nsew
rlabel metal2 s 1398 24202 1454 25002 4 i0[0]
port 3 nsew
rlabel metal2 s 4250 24202 4306 25002 4 i0[1]
port 4 nsew
rlabel metal2 s 7102 24202 7158 25002 4 i0[2]
port 5 nsew
rlabel metal2 s 9954 24202 10010 25002 4 i0[3]
port 6 nsew
rlabel metal2 s 12806 24202 12862 25002 4 i0[4]
port 7 nsew
rlabel metal2 s 15658 24202 15714 25002 4 i0[5]
port 8 nsew
rlabel metal2 s 18510 24202 18566 25002 4 i0[6]
port 9 nsew
rlabel metal2 s 21362 24202 21418 25002 4 i0[7]
port 10 nsew
rlabel metal2 s 1398 0 1454 800 4 i1[0]
port 11 nsew
rlabel metal2 s 4250 0 4306 800 4 i1[1]
port 12 nsew
rlabel metal2 s 7102 0 7158 800 4 i1[2]
port 13 nsew
rlabel metal2 s 9954 0 10010 800 4 i1[3]
port 14 nsew
rlabel metal2 s 12806 0 12862 800 4 i1[4]
port 15 nsew
rlabel metal2 s 15658 0 15714 800 4 i1[5]
port 16 nsew
rlabel metal2 s 18510 0 18566 800 4 i1[6]
port 17 nsew
rlabel metal2 s 21362 0 21418 800 4 i1[7]
port 18 nsew
rlabel metal3 s 22058 1368 22858 1488 4 s[0]
port 19 nsew
rlabel metal3 s 22058 4088 22858 4208 4 s[1]
port 20 nsew
rlabel metal3 s 22058 6808 22858 6928 4 s[2]
port 21 nsew
rlabel metal3 s 22058 9664 22858 9784 4 s[3]
port 22 nsew
rlabel metal3 s 22058 12384 22858 12504 4 s[4]
port 23 nsew
rlabel metal3 s 22058 15240 22858 15360 4 s[5]
port 24 nsew
rlabel metal3 s 22058 17960 22858 18080 4 s[6]
port 25 nsew
rlabel metal3 s 22058 20816 22858 20936 4 s[7]
port 26 nsew
rlabel metal4 s 18117 2128 18437 22352 4 VPWR
port 27 nsew
rlabel metal4 s 11248 2128 11568 22352 4 VPWR
port 27 nsew
rlabel metal4 s 4379 2128 4699 22352 4 VPWR
port 27 nsew
rlabel metal5 s 1104 18741 21712 19061 4 VPWR
port 27 nsew
rlabel metal5 s 1104 12032 21712 12352 4 VPWR
port 27 nsew
rlabel metal5 s 1104 5323 21712 5643 4 VPWR
port 27 nsew
rlabel metal4 s 14683 2128 15003 22352 4 VGND
port 28 nsew
rlabel metal4 s 7813 2128 8133 22352 4 VGND
port 28 nsew
rlabel metal5 s 1104 15387 21712 15707 4 VGND
port 28 nsew
rlabel metal5 s 1104 8677 21712 8997 4 VGND
port 28 nsew
<< properties >>
string FIXED_BBOX 0 0 22858 25002
<< end >>
