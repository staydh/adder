VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adder
  CLASS BLOCK ;
  FOREIGN adder ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.290 BY 125.010 ;
  PIN ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END ci
  PIN co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.290 117.680 114.290 118.280 ;
    END
  END co
  PIN i0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 121.010 7.270 125.010 ;
    END
  END i0[0]
  PIN i0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 121.010 21.530 125.010 ;
    END
  END i0[1]
  PIN i0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 121.010 35.790 125.010 ;
    END
  END i0[2]
  PIN i0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 121.010 50.050 125.010 ;
    END
  END i0[3]
  PIN i0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 121.010 64.310 125.010 ;
    END
  END i0[4]
  PIN i0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 121.010 78.570 125.010 ;
    END
  END i0[5]
  PIN i0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 121.010 92.830 125.010 ;
    END
  END i0[6]
  PIN i0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 121.010 107.090 125.010 ;
    END
  END i0[7]
  PIN i1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END i1[0]
  PIN i1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END i1[1]
  PIN i1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END i1[2]
  PIN i1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END i1[3]
  PIN i1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END i1[4]
  PIN i1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END i1[5]
  PIN i1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END i1[6]
  PIN i1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END i1[7]
  PIN s[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.290 6.840 114.290 7.440 ;
    END
  END s[0]
  PIN s[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.290 20.440 114.290 21.040 ;
    END
  END s[1]
  PIN s[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.290 34.040 114.290 34.640 ;
    END
  END s[2]
  PIN s[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.290 48.320 114.290 48.920 ;
    END
  END s[3]
  PIN s[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.290 61.920 114.290 62.520 ;
    END
  END s[4]
  PIN s[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.290 76.200 114.290 76.800 ;
    END
  END s[5]
  PIN s[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.290 89.800 114.290 90.400 ;
    END
  END s[6]
  PIN s[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.290 104.080 114.290 104.680 ;
    END
  END s[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 90.585 10.640 92.185 111.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 56.240 10.640 57.840 111.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.895 10.640 23.495 111.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 93.705 108.560 95.305 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 60.160 108.560 61.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.615 108.560 28.215 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.415 10.640 75.015 111.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.065 10.640 40.665 111.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 76.935 108.560 78.535 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 43.385 108.560 44.985 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 108.560 111.605 ;
      LAYER met1 ;
        RECT 5.520 4.460 108.560 111.760 ;
      LAYER met2 ;
        RECT 7.550 120.730 20.970 121.010 ;
        RECT 21.810 120.730 35.230 121.010 ;
        RECT 36.070 120.730 49.490 121.010 ;
        RECT 50.330 120.730 63.750 121.010 ;
        RECT 64.590 120.730 78.010 121.010 ;
        RECT 78.850 120.730 92.270 121.010 ;
        RECT 93.110 120.730 106.530 121.010 ;
        RECT 7.000 4.280 107.080 120.730 ;
        RECT 7.550 4.000 20.970 4.280 ;
        RECT 21.810 4.000 35.230 4.280 ;
        RECT 36.070 4.000 49.490 4.280 ;
        RECT 50.330 4.000 63.750 4.280 ;
        RECT 64.590 4.000 78.010 4.280 ;
        RECT 78.850 4.000 92.270 4.280 ;
        RECT 93.110 4.000 106.530 4.280 ;
      LAYER met3 ;
        RECT 4.000 117.280 109.890 118.145 ;
        RECT 4.000 105.080 110.290 117.280 ;
        RECT 4.000 103.680 109.890 105.080 ;
        RECT 4.000 90.800 110.290 103.680 ;
        RECT 4.000 89.400 109.890 90.800 ;
        RECT 4.000 77.200 110.290 89.400 ;
        RECT 4.000 75.800 109.890 77.200 ;
        RECT 4.000 63.600 110.290 75.800 ;
        RECT 4.400 62.920 110.290 63.600 ;
        RECT 4.400 62.200 109.890 62.920 ;
        RECT 4.000 61.520 109.890 62.200 ;
        RECT 4.000 49.320 110.290 61.520 ;
        RECT 4.000 47.920 109.890 49.320 ;
        RECT 4.000 35.040 110.290 47.920 ;
        RECT 4.000 33.640 109.890 35.040 ;
        RECT 4.000 21.440 110.290 33.640 ;
        RECT 4.000 20.040 109.890 21.440 ;
        RECT 4.000 7.840 110.290 20.040 ;
        RECT 4.000 6.975 109.890 7.840 ;
      LAYER met4 ;
        RECT 23.895 10.640 38.665 111.760 ;
        RECT 41.065 10.640 55.840 111.760 ;
        RECT 58.240 10.640 73.015 111.760 ;
      LAYER met5 ;
        RECT 5.520 63.360 108.560 75.335 ;
        RECT 5.520 46.585 108.560 58.560 ;
        RECT 5.520 29.815 108.560 41.785 ;
  END
END adder
END LIBRARY

