module adder (ci,
    co,
    VPWR,
    VGND,
    i0,
    i1,
    s);
 input ci;
 output co;
 input VPWR;
 input VGND;
 input [7:0] i0;
 input [7:0] i1;
 output [7:0] s;

 sky130_fd_sc_hd__a2bb2o_4 _25_ (.A1_N(i1[3]),
    .A2_N(i0[3]),
    .B1(i1[3]),
    .B2(i0[3]),
    .X(_00_));
 sky130_fd_sc_hd__and2_4 _26_ (.A(i0[2]),
    .B(i1[2]),
    .X(_01_));
 sky130_fd_sc_hd__and2_4 _27_ (.A(i0[1]),
    .B(i1[1]),
    .X(_02_));
 sky130_fd_sc_hd__and2_4 _28_ (.A(i0[0]),
    .B(i1[0]),
    .X(_03_));
 sky130_fd_sc_hd__o22a_4 _29_ (.A1(i0[0]),
    .A2(i1[0]),
    .B1(ci),
    .B2(_03_),
    .X(_04_));
 sky130_fd_sc_hd__o22a_4 _30_ (.A1(i0[1]),
    .A2(i1[1]),
    .B1(_02_),
    .B2(_04_),
    .X(_05_));
 sky130_fd_sc_hd__o22a_4 _31_ (.A1(i0[2]),
    .A2(i1[2]),
    .B1(_01_),
    .B2(_05_),
    .X(_06_));
 sky130_fd_sc_hd__a2bb2o_4 _32_ (.A1_N(_00_),
    .A2_N(psn_net_3),
    .B1(_00_),
    .B2(psn_net_3),
    .X(s[3]));
 sky130_fd_sc_hd__a2bb2o_4 _33_ (.A1_N(i1[4]),
    .A2_N(i0[4]),
    .B1(i1[4]),
    .B2(i0[4]),
    .X(_07_));
 sky130_fd_sc_hd__and2_4 _34_ (.A(i1[3]),
    .B(i0[3]),
    .X(_08_));
 sky130_fd_sc_hd__o22a_4 _35_ (.A1(i1[3]),
    .A2(i0[3]),
    .B1(_08_),
    .B2(_06_),
    .X(_09_));
 sky130_fd_sc_hd__a2bb2o_4 _36_ (.A1_N(_07_),
    .A2_N(psn_net_2),
    .B1(_07_),
    .B2(psn_net_2),
    .X(s[4]));
 sky130_fd_sc_hd__a2bb2o_4 _37_ (.A1_N(i1[5]),
    .A2_N(i0[5]),
    .B1(i1[5]),
    .B2(i0[5]),
    .X(_10_));
 sky130_fd_sc_hd__and2_4 _38_ (.A(i1[4]),
    .B(i0[4]),
    .X(_11_));
 sky130_fd_sc_hd__o22a_4 _39_ (.A1(i1[4]),
    .A2(i0[4]),
    .B1(_11_),
    .B2(_09_),
    .X(_12_));
 sky130_fd_sc_hd__a2bb2o_4 _40_ (.A1_N(_10_),
    .A2_N(psn_net_1),
    .B1(_10_),
    .B2(psn_net_1),
    .X(s[5]));
 sky130_fd_sc_hd__a2bb2o_4 _41_ (.A1_N(i1[6]),
    .A2_N(i0[6]),
    .B1(i1[6]),
    .B2(i0[6]),
    .X(_13_));
 sky130_fd_sc_hd__and2_4 _42_ (.A(i1[5]),
    .B(i0[5]),
    .X(_14_));
 sky130_fd_sc_hd__o22a_4 _43_ (.A1(i1[5]),
    .A2(i0[5]),
    .B1(_14_),
    .B2(_12_),
    .X(_15_));
 sky130_fd_sc_hd__a2bb2o_4 _44_ (.A1_N(_13_),
    .A2_N(psn_net_0),
    .B1(_13_),
    .B2(psn_net_0),
    .X(s[6]));
 sky130_fd_sc_hd__and2_4 _45_ (.A(i0[7]),
    .B(i1[7]),
    .X(_16_));
 sky130_fd_sc_hd__and2_4 _46_ (.A(i1[6]),
    .B(i0[6]),
    .X(_17_));
 sky130_fd_sc_hd__o22a_4 _47_ (.A1(i1[6]),
    .A2(i0[6]),
    .B1(_17_),
    .B2(_15_),
    .X(_18_));
 sky130_fd_sc_hd__o22a_4 _48_ (.A1(i0[7]),
    .A2(i1[7]),
    .B1(_16_),
    .B2(_18_),
    .X(co));
 sky130_fd_sc_hd__a2bb2o_4 _49_ (.A1_N(i0[7]),
    .A2_N(i1[7]),
    .B1(i0[7]),
    .B2(i1[7]),
    .X(_19_));
 sky130_fd_sc_hd__a2bb2o_4 _50_ (.A1_N(_19_),
    .A2_N(_18_),
    .B1(_18_),
    .B2(_19_),
    .X(s[7]));
 sky130_fd_sc_hd__inv_2 _51_ (.A(ci),
    .Y(_20_));
 sky130_fd_sc_hd__inv_2 _52_ (.A(psn_net_6),
    .Y(_21_));
 sky130_fd_sc_hd__o21a_4 _53_ (.A1(i0[0]),
    .A2(i1[0]),
    .B1(_21_),
    .X(_22_));
 sky130_fd_sc_hd__a2bb2o_4 _54_ (.A1_N(_20_),
    .A2_N(_22_),
    .B1(_20_),
    .B2(_22_),
    .X(s[0]));
 sky130_fd_sc_hd__a2bb2o_4 _55_ (.A1_N(i0[1]),
    .A2_N(i1[1]),
    .B1(i0[1]),
    .B2(i1[1]),
    .X(_23_));
 sky130_fd_sc_hd__a2bb2o_4 _56_ (.A1_N(_23_),
    .A2_N(psn_net_5),
    .B1(psn_net_5),
    .B2(_23_),
    .X(s[1]));
 sky130_fd_sc_hd__a2bb2o_4 _57_ (.A1_N(i0[2]),
    .A2_N(i1[2]),
    .B1(i0[2]),
    .B2(i1[2]),
    .X(_24_));
 sky130_fd_sc_hd__a2bb2o_4 _58_ (.A1_N(_24_),
    .A2_N(psn_net_4),
    .B1(psn_net_4),
    .B2(_24_),
    .X(s[2]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_209 ();
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_0 (.A(_15_),
    .X(psn_net_0));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_1 (.A(psn_net_7),
    .X(psn_net_1));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_2 (.A(psn_net_8),
    .X(psn_net_2));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_3 (.A(psn_net_9),
    .X(psn_net_3));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_4 (.A(psn_net_10),
    .X(psn_net_4));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_5 (.A(psn_net_11),
    .X(psn_net_5));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_6 (.A(psn_net_12),
    .X(psn_net_6));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_7 (.A(psn_net_13),
    .X(psn_net_7));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_8 (.A(psn_net_14),
    .X(psn_net_8));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_9 (.A(psn_net_15),
    .X(psn_net_9));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_10 (.A(psn_net_16),
    .X(psn_net_10));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_11 (.A(psn_net_17),
    .X(psn_net_11));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_12 (.A(psn_net_18),
    .X(psn_net_12));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_13 (.A(_12_),
    .X(psn_net_13));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_14 (.A(psn_net_19),
    .X(psn_net_14));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_15 (.A(psn_net_20),
    .X(psn_net_15));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_16 (.A(psn_net_21),
    .X(psn_net_16));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_17 (.A(psn_net_22),
    .X(psn_net_17));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_18 (.A(psn_net_23),
    .X(psn_net_18));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_19 (.A(psn_net_24),
    .X(psn_net_19));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_20 (.A(psn_net_25),
    .X(psn_net_20));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_21 (.A(psn_net_26),
    .X(psn_net_21));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_22 (.A(psn_net_27),
    .X(psn_net_22));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_23 (.A(psn_net_28),
    .X(psn_net_23));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_24 (.A(_09_),
    .X(psn_net_24));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_25 (.A(psn_net_29),
    .X(psn_net_25));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_26 (.A(psn_net_30),
    .X(psn_net_26));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_27 (.A(psn_net_31),
    .X(psn_net_27));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_28 (.A(psn_net_32),
    .X(psn_net_28));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_29 (.A(_06_),
    .X(psn_net_29));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_30 (.A(psn_net_33),
    .X(psn_net_30));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_31 (.A(psn_net_34),
    .X(psn_net_31));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_32 (.A(psn_net_35),
    .X(psn_net_32));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_33 (.A(_05_),
    .X(psn_net_33));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_34 (.A(psn_net_36),
    .X(psn_net_34));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_35 (.A(psn_net_37),
    .X(psn_net_35));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_36 (.A(_04_),
    .X(psn_net_36));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_37 (.A(psn_net_38),
    .X(psn_net_37));
 sky130_fd_sc_hd__buf_2 psn_inst_psn_buff_38 (.A(_03_),
    .X(psn_net_38));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_94 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_187 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_60 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_67 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_91 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_25 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_49 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_78 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_90 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_114 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_220 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_91 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_26 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_77 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_89 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_121 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_87 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_119 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_11 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_75 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_99 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_118 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_220 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_108 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_120 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_152 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_119 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_220 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_119 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_151 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_90 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_121 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_220 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_106 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_130 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_149 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_131 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_220 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_150 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_150 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_182 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_220 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_151 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_178 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_136 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_148 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_220 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_162 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_181 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_179 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_220 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_185 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_155 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_182 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_220 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_162 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_213 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_218 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_192 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_220 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_213 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_44 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_68 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_80 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_93 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_105 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_129 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_154 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_166 ();
 sky130_fd_sc_hd__decap_12 FILLER_34_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_215 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_62 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_74 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_86 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_123 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_147 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_159 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_35_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_213 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_32 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_63 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_87 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_94 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_118 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_125 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_149 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_180 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_187 ();
 sky130_fd_sc_hd__decap_12 FILLER_36_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_218 ();
endmodule
