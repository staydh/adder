magic
tech sky130A
magscale 1 2
timestamp 1616762078
<< obsli1 >>
rect 1104 2159 21712 22321
<< obsm1 >>
rect 1104 892 21712 22352
<< metal2 >>
rect 1398 24202 1454 25002
rect 4250 24202 4306 25002
rect 7102 24202 7158 25002
rect 9954 24202 10010 25002
rect 12806 24202 12862 25002
rect 15658 24202 15714 25002
rect 18510 24202 18566 25002
rect 21362 24202 21418 25002
rect 1398 0 1454 800
rect 4250 0 4306 800
rect 7102 0 7158 800
rect 9954 0 10010 800
rect 12806 0 12862 800
rect 15658 0 15714 800
rect 18510 0 18566 800
rect 21362 0 21418 800
<< obsm2 >>
rect 1510 24146 4194 24202
rect 4362 24146 7046 24202
rect 7214 24146 9898 24202
rect 10066 24146 12750 24202
rect 12918 24146 15602 24202
rect 15770 24146 18454 24202
rect 18622 24146 21306 24202
rect 1400 856 21416 24146
rect 1510 800 4194 856
rect 4362 800 7046 856
rect 7214 800 9898 856
rect 10066 800 12750 856
rect 12918 800 15602 856
rect 15770 800 18454 856
rect 18622 800 21306 856
<< metal3 >>
rect 22058 23536 22858 23656
rect 22058 20816 22858 20936
rect 22058 17960 22858 18080
rect 22058 15240 22858 15360
rect 0 12520 800 12640
rect 22058 12384 22858 12504
rect 22058 9664 22858 9784
rect 22058 6808 22858 6928
rect 22058 4088 22858 4208
rect 22058 1368 22858 1488
<< obsm3 >>
rect 800 23456 21978 23629
rect 800 21016 22058 23456
rect 800 20736 21978 21016
rect 800 18160 22058 20736
rect 800 17880 21978 18160
rect 800 15440 22058 17880
rect 800 15160 21978 15440
rect 800 12720 22058 15160
rect 880 12584 22058 12720
rect 880 12440 21978 12584
rect 800 12304 21978 12440
rect 800 9864 22058 12304
rect 800 9584 21978 9864
rect 800 7008 22058 9584
rect 800 6728 21978 7008
rect 800 4288 22058 6728
rect 800 4008 21978 4288
rect 800 1568 22058 4008
rect 800 1395 21978 1568
<< metal4 >>
rect 4379 2128 4699 22352
rect 7813 2128 8133 22352
rect 11248 2128 11568 22352
rect 14683 2128 15003 22352
rect 18117 2128 18437 22352
<< obsm4 >>
rect 4779 2128 7733 22352
rect 8213 2128 11168 22352
rect 11648 2128 14603 22352
<< metal5 >>
rect 1104 18741 21712 19061
rect 1104 15387 21712 15707
rect 1104 12032 21712 12352
rect 1104 8677 21712 8997
rect 1104 5323 21712 5643
<< obsm5 >>
rect 1104 12672 21712 15067
rect 1104 9317 21712 11712
rect 1104 5963 21712 8357
<< labels >>
rlabel metal3 s 0 12520 800 12640 6 ci
port 1 nsew signal input
rlabel metal3 s 22058 23536 22858 23656 6 co
port 2 nsew signal output
rlabel metal2 s 1398 24202 1454 25002 6 i0[0]
port 3 nsew signal input
rlabel metal2 s 4250 24202 4306 25002 6 i0[1]
port 4 nsew signal input
rlabel metal2 s 7102 24202 7158 25002 6 i0[2]
port 5 nsew signal input
rlabel metal2 s 9954 24202 10010 25002 6 i0[3]
port 6 nsew signal input
rlabel metal2 s 12806 24202 12862 25002 6 i0[4]
port 7 nsew signal input
rlabel metal2 s 15658 24202 15714 25002 6 i0[5]
port 8 nsew signal input
rlabel metal2 s 18510 24202 18566 25002 6 i0[6]
port 9 nsew signal input
rlabel metal2 s 21362 24202 21418 25002 6 i0[7]
port 10 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 i1[0]
port 11 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 i1[1]
port 12 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 i1[2]
port 13 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 i1[3]
port 14 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 i1[4]
port 15 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 i1[5]
port 16 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 i1[6]
port 17 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 i1[7]
port 18 nsew signal input
rlabel metal3 s 22058 1368 22858 1488 6 s[0]
port 19 nsew signal output
rlabel metal3 s 22058 4088 22858 4208 6 s[1]
port 20 nsew signal output
rlabel metal3 s 22058 6808 22858 6928 6 s[2]
port 21 nsew signal output
rlabel metal3 s 22058 9664 22858 9784 6 s[3]
port 22 nsew signal output
rlabel metal3 s 22058 12384 22858 12504 6 s[4]
port 23 nsew signal output
rlabel metal3 s 22058 15240 22858 15360 6 s[5]
port 24 nsew signal output
rlabel metal3 s 22058 17960 22858 18080 6 s[6]
port 25 nsew signal output
rlabel metal3 s 22058 20816 22858 20936 6 s[7]
port 26 nsew signal output
rlabel metal4 s 18117 2128 18437 22352 6 VPWR
port 27 nsew power bidirectional
rlabel metal4 s 11248 2128 11568 22352 6 VPWR
port 28 nsew power bidirectional
rlabel metal4 s 4379 2128 4699 22352 6 VPWR
port 29 nsew power bidirectional
rlabel metal5 s 1104 18741 21712 19061 6 VPWR
port 30 nsew power bidirectional
rlabel metal5 s 1104 12032 21712 12352 6 VPWR
port 31 nsew power bidirectional
rlabel metal5 s 1104 5323 21712 5643 6 VPWR
port 32 nsew power bidirectional
rlabel metal4 s 14683 2128 15003 22352 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 7813 2128 8133 22352 6 VGND
port 34 nsew ground bidirectional
rlabel metal5 s 1104 15387 21712 15707 6 VGND
port 35 nsew ground bidirectional
rlabel metal5 s 1104 8677 21712 8997 6 VGND
port 36 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 22858 25002
string LEFview TRUE
<< end >>
