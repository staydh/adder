# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

# High density, single height
SITE unithd
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 2.72 ;
END unithd

# High density, double height
SITE unithddbl
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.46 0.34 ;
  OFFSET 0.23 0.17 ;

  WIDTH 0.17 ;          # LI 1
  # SPACING  0.17 ;     # LI 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.17 ;
  AREA 0.0561 ;         # LI 6
  THICKNESS 0.1 ;
  EDGECAPACITANCE 40.697E-6 ;
  CAPACITANCE CPERSQDIST 36.9866E-6 ;
  RESISTANCE RPERSQ 12.2 ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 75 ) ( 0.0125 75 ) ( 0.0225 85.125 ) ( 22.5 10200 ) ) ;
END li1

LAYER mcon
  TYPE CUT ;

  WIDTH 0.17 ;                # Mcon 1
  SPACING 0.19 ;              # Mcon 2
  ENCLOSURE BELOW 0 0 ;       # Mcon 4
  ENCLOSURE ABOVE 0.03 0.06 ; # Met1 4 / Met1 5

  ANTENNADIFFAREARATIO PWL ( ( 0 3 ) ( 0.0125 3 ) ( 0.0225 3.405 ) ( 22.5 408 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.36 ; # mA per via Iavg_max at Tj = 90oC

END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.34 ;
  OFFSET 0.17 ;

  WIDTH 0.14 ;                     # Met1 1
  # SPACING 0.14 ;                 # Met1 2
  # SPACING 0.28 RANGE 3.001 100 ; # Met1 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.083 ;                     # Met1 6
  THICKNESS 0.35 ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  EDGECAPACITANCE 40.567E-6 ;
  CAPACITANCE CPERSQDIST 25.7784E-6 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;

  RESISTANCE RPERSQ 0.125 ;
END met1

LAYER via
  TYPE CUT ;
  WIDTH 0.15 ;                  # Via 1a
  SPACING 0.17 ;                # Via 2
  ENCLOSURE BELOW 0.055 0.085 ; # Via 4a / Via 5a
  ENCLOSURE ABOVE 0.055 0.085 ; # Met2 4 / Met2 5

  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.29 ; # mA per via Iavg_max at Tj = 90oC
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.46 ;
  OFFSET 0.23 ;

  WIDTH 0.14 ;                        # Met2 1
  # SPACING  0.14 ;                   # Met2 2
  # SPACING  0.28 RANGE 3.001 100 ;   # Met2 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.0676 ;                       # Met2 6
  THICKNESS 0.35 ;

  EDGECAPACITANCE 37.759E-6 ;
  CAPACITANCE CPERSQDIST 16.9423E-6 ;
  RESISTANCE RPERSQ 0.125 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met2

# ******** Layer via2, type routing, number 44 **************
LAYER via2
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via2 1
  SPACING 0.2 ;                 # Via2 2
  ENCLOSURE BELOW 0.04 0.085 ;  # Via2 4
  ENCLOSURE ABOVE 0.065 0.065 ; # Met3 4
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.68 ;
  OFFSET 0.34 ;

  WIDTH 0.3 ;              # Met3 1
  # SPACING 0.3 ;          # Met3 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;              # Met3 6
  THICKNESS 0.8 ;

  EDGECAPACITANCE 40.989E-6 ;
  CAPACITANCE CPERSQDIST 12.3729E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met3

LAYER via3
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via3 1
  SPACING 0.2 ;                 # Via3 2
  ENCLOSURE BELOW 0.06 0.09 ;   # Via3 4 / Via3 5
  ENCLOSURE ABOVE 0.065 0.065 ; # Met4 3
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.92 ;
  OFFSET 0.46 ;

  WIDTH 0.3 ;             # Met4 1
  # SPACING  0.3 ;             # Met4 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;            # Met4 4a

  THICKNESS 0.8 ;

  EDGECAPACITANCE 36.676E-6 ;
  CAPACITANCE CPERSQDIST 8.41537E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met4

LAYER via4
  TYPE CUT ;

  WIDTH 0.8 ;                 # Via4 1
  SPACING 0.8 ;               # Via4 2
  ENCLOSURE BELOW 0.19 0.19 ; # Via4 4
  ENCLOSURE ABOVE 0.31 0.31 ; # Met5 3
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 2.49 ; # mA per via Iavg_max at Tj = 90oC
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 3.4 ;
  OFFSET 1.7 ;

  WIDTH 1.6 ;            # Met5 1
  #SPACING  1.6 ;        # Met5 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 1.6 ;
  AREA 4 ;               # Met5 4

  THICKNESS 1.2 ;

  EDGECAPACITANCE 38.851E-6 ;
  CAPACITANCE CPERSQDIST 6.32063E-6 ;
  RESISTANCE RPERSQ 0.0285 ;
  DCCURRENTDENSITY AVERAGE 10.17 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 22.34 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met5


### Routing via cells section   ###
# Plus via rule, metals are along the prefered direction
VIA L1M1_PR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIARULE L1M1_PR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR

# Plus via rule, metals are along the non prefered direction
VIA L1M1_PR_R DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIARULE L1M1_PR_R GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA L1M1_PR_M DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIARULE L1M1_PR_M GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA L1M1_PR_MR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIARULE L1M1_PR_MR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_MR

# Centered via rule, we really do not want to use it
VIA L1M1_PR_C DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIARULE L1M1_PR_C GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_C

# Plus via rule, metals are along the prefered direction
VIA M1M2_PR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIARULE M1M2_PR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR

# Plus via rule, metals are along the non prefered direction
VIA M1M2_PR_R DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIARULE M1M2_PR_R GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M1M2_PR_M DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIARULE M1M2_PR_M GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M1M2_PR_MR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIARULE M1M2_PR_MR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_MR

# Centered via rule, we really do not want to use it
VIA M1M2_PR_C DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.16 0.16 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIARULE M1M2_PR_C GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_C

# Plus via rule, metals are along the prefered direction
VIA M2M3_PR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIARULE M2M3_PR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR

# Plus via rule, metals are along the non prefered direction
VIA M2M3_PR_R DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIARULE M2M3_PR_R GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M2M3_PR_M DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIARULE M2M3_PR_M GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M2M3_PR_MR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIARULE M2M3_PR_MR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_MR

# Centered via rule, we really do not want to use it
VIA M2M3_PR_C DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.185 0.185 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIARULE M2M3_PR_C GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_C

# Plus via rule, metals are along the prefered direction
VIA M3M4_PR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIARULE M3M4_PR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR

# Plus via rule, metals are along the non prefered direction
VIA M3M4_PR_R DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIARULE M3M4_PR_R GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M3M4_PR_M DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIARULE M3M4_PR_M GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M3M4_PR_MR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIARULE M3M4_PR_MR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_MR

# Centered via rule, we really do not want to use it
VIA M3M4_PR_C DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.19 0.19 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIARULE M3M4_PR_C GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_C

# Plus via rule, metals are along the prefered direction
VIA M4M5_PR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIARULE M4M5_PR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR

# Plus via rule, metals are along the non prefered direction
VIA M4M5_PR_R DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIARULE M4M5_PR_R GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M4M5_PR_M DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIARULE M4M5_PR_M GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M4M5_PR_MR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIARULE M4M5_PR_MR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_MR

# Centered via rule, we really do not want to use it
VIA M4M5_PR_C DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

VIARULE M4M5_PR_C GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_C
###  end of single via cells   ###


MACRO sky130_ef_sc_hd__fakediode_2
  CLASS CORE SPACER ;
  FOREIGN sky130_ef_sc_hd__fakediode_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIODE
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.835 2.465 ;
    END
  END DIODE
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.920 0.085 ;
      LAYER mcon ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.920 0.240 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 0.920 2.805 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.960 ;
    END
  END VPWR
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.110 2.910 ;
    END
  END VPB
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
END sky130_ef_sc_hd__fakediode_2
MACRO sky130_fd_sc_hd__sdfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.34000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.575000 0.265000 11.925000 1.695000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.435000 1.535000 12.825000 2.080000 ;
        RECT 12.445000 0.310000 12.825000 0.825000 ;
        RECT 12.525000 2.080000 12.825000 2.465000 ;
        RECT 12.655000 0.825000 12.825000 1.535000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
      LAYER mcon ;
        RECT 6.865000 0.765000 7.035000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
      LAYER mcon ;
        RECT 9.690000 1.105000  9.860000 1.275000 ;
        RECT 9.945000 0.765000 10.115000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215000 -0.010000 0.235000 0.015000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  1.970000 1.425000 ;
        RECT -0.190000 1.425000 13.530000 2.910000 ;
        RECT  4.405000 1.305000 13.530000 1.425000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.340000 0.085000 ;
      RECT  0.000000  2.635000 13.340000 2.805000 ;
      RECT  0.090000  1.795000  0.865000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.530000  2.135000  0.860000 2.635000 ;
      RECT  0.660000  0.805000  0.835000 0.995000 ;
      RECT  0.660000  0.995000  0.975000 1.325000 ;
      RECT  0.660000  1.325000  0.865000 1.795000 ;
      RECT  1.015000  0.345000  1.315000 0.675000 ;
      RECT  1.035000  1.730000  1.315000 1.900000 ;
      RECT  1.035000  1.900000  1.205000 2.465000 ;
      RECT  1.145000  0.675000  1.315000 1.730000 ;
      RECT  1.535000  0.395000  1.705000 0.730000 ;
      RECT  1.535000  0.730000  2.225000 0.900000 ;
      RECT  1.875000  0.085000  2.205000 0.560000 ;
      RECT  1.900000  2.055000  2.150000 2.400000 ;
      RECT  1.980000  1.260000  2.470000 1.455000 ;
      RECT  1.980000  1.455000  2.150000 2.055000 ;
      RECT  2.055000  0.900000  2.225000 0.995000 ;
      RECT  2.055000  0.995000  3.085000 1.185000 ;
      RECT  2.055000  1.185000  2.470000 1.260000 ;
      RECT  2.320000  2.040000  2.490000 2.635000 ;
      RECT  2.395000  0.085000  2.725000 0.825000 ;
      RECT  2.915000  0.255000  3.850000 0.425000 ;
      RECT  2.915000  0.425000  3.085000 0.995000 ;
      RECT  3.255000  0.675000  3.425000 1.015000 ;
      RECT  3.255000  1.015000  3.460000 1.185000 ;
      RECT  3.290000  1.185000  3.460000 1.935000 ;
      RECT  3.290000  1.935000  5.075000 2.105000 ;
      RECT  3.460000  2.105000  3.630000 2.465000 ;
      RECT  3.680000  0.425000  3.850000 1.685000 ;
      RECT  4.300000  2.275000  4.630000 2.635000 ;
      RECT  4.445000  0.085000  4.775000 0.540000 ;
      RECT  4.565000  0.715000  5.145000 0.895000 ;
      RECT  4.565000  0.895000  4.735000 1.935000 ;
      RECT  4.905000  1.065000  5.075000 1.395000 ;
      RECT  4.905000  2.105000  5.075000 2.185000 ;
      RECT  4.905000  2.185000  5.275000 2.435000 ;
      RECT  4.975000  0.335000  5.315000 0.505000 ;
      RECT  4.975000  0.505000  5.145000 0.715000 ;
      RECT  5.245000  1.575000  5.495000 1.955000 ;
      RECT  5.325000  0.705000  5.975000 1.035000 ;
      RECT  5.325000  1.035000  5.495000 1.575000 ;
      RECT  5.470000  2.135000  5.835000 2.465000 ;
      RECT  5.485000  0.305000  6.335000 0.475000 ;
      RECT  5.665000  1.215000  7.375000 1.385000 ;
      RECT  5.665000  1.385000  5.835000 2.135000 ;
      RECT  6.005000  1.935000  7.165000 2.105000 ;
      RECT  6.005000  2.105000  6.175000 2.375000 ;
      RECT  6.165000  0.475000  6.335000 1.215000 ;
      RECT  6.285000  1.595000  7.715000 1.765000 ;
      RECT  6.410000  2.355000  6.740000 2.635000 ;
      RECT  6.915000  0.085000  7.245000 0.545000 ;
      RECT  6.995000  2.105000  7.165000 2.375000 ;
      RECT  7.205000  1.005000  7.375000 1.215000 ;
      RECT  7.375000  2.175000  7.745000 2.635000 ;
      RECT  7.455000  0.275000  7.785000 0.445000 ;
      RECT  7.455000  0.445000  7.715000 0.835000 ;
      RECT  7.455000  1.765000  7.715000 1.835000 ;
      RECT  7.455000  1.835000  8.140000 2.005000 ;
      RECT  7.545000  0.835000  7.715000 1.595000 ;
      RECT  7.885000  0.705000  8.095000 1.495000 ;
      RECT  7.885000  1.495000  8.520000 1.655000 ;
      RECT  7.885000  1.655000  8.870000 1.665000 ;
      RECT  7.970000  2.005000  8.140000 2.465000 ;
      RECT  8.005000  0.255000  8.915000 0.535000 ;
      RECT  8.310000  1.665000  8.870000 1.935000 ;
      RECT  8.310000  1.935000  8.840000 1.955000 ;
      RECT  8.320000  2.125000  9.190000 2.465000 ;
      RECT  8.405000  0.920000  8.575000 1.325000 ;
      RECT  8.745000  0.535000  8.915000 1.315000 ;
      RECT  8.745000  1.315000  9.210000 1.485000 ;
      RECT  9.015000  2.035000  9.210000 2.115000 ;
      RECT  9.015000  2.115000  9.190000 2.125000 ;
      RECT  9.040000  1.485000  9.210000 1.575000 ;
      RECT  9.040000  1.575000 10.205000 1.745000 ;
      RECT  9.040000  1.745000  9.210000 2.035000 ;
      RECT  9.085000  0.085000  9.255000 0.525000 ;
      RECT  9.125000  0.695000  9.655000 0.865000 ;
      RECT  9.125000  0.865000  9.295000 1.145000 ;
      RECT  9.360000  2.195000  9.610000 2.635000 ;
      RECT  9.485000  0.295000 10.515000 0.465000 ;
      RECT  9.485000  0.465000  9.655000 0.695000 ;
      RECT  9.780000  1.915000 10.545000 2.085000 ;
      RECT  9.780000  2.085000  9.950000 2.375000 ;
      RECT 10.120000  2.255000 10.450000 2.635000 ;
      RECT 10.345000  0.465000 10.515000 1.055000 ;
      RECT 10.345000  1.055000 11.060000 1.295000 ;
      RECT 10.375000  1.295000 11.060000 1.325000 ;
      RECT 10.375000  1.325000 10.545000 1.915000 ;
      RECT 10.715000  0.345000 10.885000 0.715000 ;
      RECT 10.715000  0.715000 11.405000 0.885000 ;
      RECT 10.715000  1.795000 11.405000 1.865000 ;
      RECT 10.715000  1.865000 12.265000 2.035000 ;
      RECT 10.715000  2.035000 10.890000 2.465000 ;
      RECT 11.090000  0.085000 11.365000 0.545000 ;
      RECT 11.090000  2.205000 11.420000 2.635000 ;
      RECT 11.230000  0.885000 11.405000 1.795000 ;
      RECT 11.550000  2.035000 12.265000 2.085000 ;
      RECT 12.025000  2.255000 12.355000 2.635000 ;
      RECT 12.095000  0.995000 12.485000 1.325000 ;
      RECT 12.095000  1.325000 12.265000 1.865000 ;
      RECT 12.105000  0.085000 12.275000 0.825000 ;
      RECT 12.995000  0.085000 13.165000 0.930000 ;
      RECT 12.995000  1.495000 13.245000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.805000  1.105000  0.975000 1.275000 ;
      RECT  1.035000  1.785000  1.205000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.905000  1.105000  5.075000 1.275000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.325000  1.785000  5.495000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.405000  1.105000  8.575000 1.275000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.445000  1.785000  8.615000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
    LAYER met1 ;
      RECT 0.745000 1.075000 1.035000 1.120000 ;
      RECT 0.745000 1.120000 8.635000 1.260000 ;
      RECT 0.745000 1.260000 1.035000 1.305000 ;
      RECT 0.970000 1.755000 1.270000 1.800000 ;
      RECT 0.970000 1.800000 8.675000 1.940000 ;
      RECT 0.970000 1.940000 1.270000 1.985000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrbp_2
MACRO sky130_fd_sc_hd__sdfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.88000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.140000 0.265000 11.400000 0.795000 ;
        RECT 11.140000 1.460000 11.400000 2.325000 ;
        RECT 11.150000 1.445000 11.400000 1.460000 ;
        RECT 11.190000 0.795000 11.400000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.510000 1.560000 12.780000 2.465000 ;
        RECT 12.520000 0.255000 12.780000 0.760000 ;
        RECT 12.600000 0.760000 12.780000 1.560000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
      LAYER mcon ;
        RECT 6.865000 0.765000 7.035000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
      LAYER mcon ;
        RECT 9.690000 1.105000  9.860000 1.275000 ;
        RECT 9.945000 0.765000 10.115000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215000 -0.010000 0.235000 0.015000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  1.970000 1.425000 ;
        RECT -0.190000 1.425000 13.070000 2.910000 ;
        RECT  4.405000 1.305000 13.070000 1.425000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.880000 0.085000 ;
      RECT  0.000000  2.635000 12.880000 2.805000 ;
      RECT  0.090000  1.795000  0.865000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.530000  2.135000  0.860000 2.635000 ;
      RECT  0.660000  0.805000  0.835000 0.995000 ;
      RECT  0.660000  0.995000  0.975000 1.325000 ;
      RECT  0.660000  1.325000  0.865000 1.795000 ;
      RECT  1.015000  0.345000  1.315000 0.675000 ;
      RECT  1.035000  1.730000  1.315000 1.900000 ;
      RECT  1.035000  1.900000  1.205000 2.465000 ;
      RECT  1.145000  0.675000  1.315000 1.730000 ;
      RECT  1.535000  0.395000  1.705000 0.730000 ;
      RECT  1.535000  0.730000  2.225000 0.900000 ;
      RECT  1.875000  0.085000  2.205000 0.560000 ;
      RECT  1.900000  2.055000  2.150000 2.400000 ;
      RECT  1.980000  1.260000  2.470000 1.455000 ;
      RECT  1.980000  1.455000  2.150000 2.055000 ;
      RECT  2.055000  0.900000  2.225000 0.995000 ;
      RECT  2.055000  0.995000  3.085000 1.185000 ;
      RECT  2.055000  1.185000  2.470000 1.260000 ;
      RECT  2.320000  2.040000  2.490000 2.635000 ;
      RECT  2.395000  0.085000  2.725000 0.825000 ;
      RECT  2.915000  0.255000  3.850000 0.425000 ;
      RECT  2.915000  0.425000  3.085000 0.995000 ;
      RECT  3.255000  0.675000  3.425000 1.015000 ;
      RECT  3.255000  1.015000  3.460000 1.185000 ;
      RECT  3.290000  1.185000  3.460000 1.935000 ;
      RECT  3.290000  1.935000  5.075000 2.105000 ;
      RECT  3.460000  2.105000  3.630000 2.465000 ;
      RECT  3.680000  0.425000  3.850000 1.685000 ;
      RECT  4.300000  2.275000  4.630000 2.635000 ;
      RECT  4.445000  0.085000  4.775000 0.540000 ;
      RECT  4.565000  0.715000  5.145000 0.895000 ;
      RECT  4.565000  0.895000  4.735000 1.935000 ;
      RECT  4.905000  1.065000  5.075000 1.395000 ;
      RECT  4.905000  2.105000  5.075000 2.185000 ;
      RECT  4.905000  2.185000  5.275000 2.435000 ;
      RECT  4.975000  0.335000  5.315000 0.505000 ;
      RECT  4.975000  0.505000  5.145000 0.715000 ;
      RECT  5.245000  1.575000  5.495000 1.955000 ;
      RECT  5.325000  0.705000  5.975000 1.035000 ;
      RECT  5.325000  1.035000  5.495000 1.575000 ;
      RECT  5.470000  2.135000  5.835000 2.465000 ;
      RECT  5.485000  0.305000  6.335000 0.475000 ;
      RECT  5.665000  1.215000  7.375000 1.385000 ;
      RECT  5.665000  1.385000  5.835000 2.135000 ;
      RECT  6.005000  1.935000  7.165000 2.105000 ;
      RECT  6.005000  2.105000  6.175000 2.375000 ;
      RECT  6.165000  0.475000  6.335000 1.215000 ;
      RECT  6.285000  1.595000  7.715000 1.765000 ;
      RECT  6.410000  2.355000  6.740000 2.635000 ;
      RECT  6.915000  0.085000  7.245000 0.545000 ;
      RECT  6.995000  2.105000  7.165000 2.375000 ;
      RECT  7.205000  1.005000  7.375000 1.215000 ;
      RECT  7.375000  2.175000  7.745000 2.635000 ;
      RECT  7.455000  0.275000  7.785000 0.445000 ;
      RECT  7.455000  0.445000  7.715000 0.835000 ;
      RECT  7.455000  1.765000  7.715000 1.835000 ;
      RECT  7.455000  1.835000  8.140000 2.005000 ;
      RECT  7.545000  0.835000  7.715000 1.595000 ;
      RECT  7.885000  0.705000  8.095000 1.495000 ;
      RECT  7.885000  1.495000  8.520000 1.655000 ;
      RECT  7.885000  1.655000  8.870000 1.665000 ;
      RECT  7.970000  2.005000  8.140000 2.465000 ;
      RECT  8.005000  0.255000  8.915000 0.535000 ;
      RECT  8.310000  1.665000  8.870000 1.935000 ;
      RECT  8.310000  1.935000  8.840000 1.955000 ;
      RECT  8.320000  2.125000  9.190000 2.465000 ;
      RECT  8.405000  0.920000  8.575000 1.325000 ;
      RECT  8.745000  0.535000  8.915000 1.315000 ;
      RECT  8.745000  1.315000  9.210000 1.485000 ;
      RECT  9.015000  2.035000  9.210000 2.115000 ;
      RECT  9.015000  2.115000  9.190000 2.125000 ;
      RECT  9.040000  1.485000  9.210000 1.575000 ;
      RECT  9.040000  1.575000 10.205000 1.745000 ;
      RECT  9.040000  1.745000  9.210000 2.035000 ;
      RECT  9.085000  0.085000  9.255000 0.525000 ;
      RECT  9.125000  0.695000  9.655000 0.865000 ;
      RECT  9.125000  0.865000  9.295000 1.145000 ;
      RECT  9.360000  2.195000  9.610000 2.635000 ;
      RECT  9.485000  0.295000 10.515000 0.465000 ;
      RECT  9.485000  0.465000  9.655000 0.695000 ;
      RECT  9.780000  1.915000 10.545000 2.085000 ;
      RECT  9.780000  2.085000  9.950000 2.375000 ;
      RECT 10.120000  2.255000 10.450000 2.635000 ;
      RECT 10.345000  0.465000 10.515000 0.995000 ;
      RECT 10.345000  0.995000 11.020000 1.295000 ;
      RECT 10.375000  1.295000 11.020000 1.325000 ;
      RECT 10.375000  1.325000 10.545000 1.915000 ;
      RECT 10.720000  0.085000 10.890000 0.545000 ;
      RECT 10.720000  1.495000 10.970000 2.635000 ;
      RECT 11.650000  1.535000 12.325000 1.705000 ;
      RECT 11.650000  1.705000 11.830000 2.465000 ;
      RECT 11.660000  0.255000 11.830000 0.635000 ;
      RECT 11.660000  0.635000 12.325000 0.805000 ;
      RECT 12.010000  0.085000 12.340000 0.465000 ;
      RECT 12.010000  1.875000 12.340000 2.635000 ;
      RECT 12.155000  0.805000 12.325000 1.060000 ;
      RECT 12.155000  1.060000 12.430000 1.390000 ;
      RECT 12.155000  1.390000 12.325000 1.535000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.805000  1.105000  0.975000 1.275000 ;
      RECT  1.035000  1.785000  1.205000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.905000  1.105000  5.075000 1.275000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.325000  1.785000  5.495000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.405000  1.105000  8.575000 1.275000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.445000  1.785000  8.615000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
    LAYER met1 ;
      RECT 0.745000 1.075000 1.035000 1.120000 ;
      RECT 0.745000 1.120000 8.635000 1.260000 ;
      RECT 0.745000 1.260000 1.035000 1.305000 ;
      RECT 0.970000 1.755000 1.270000 1.800000 ;
      RECT 0.970000 1.800000 8.675000 1.940000 ;
      RECT 0.970000 1.940000 1.270000 1.985000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrbp_1
MACRO sky130_fd_sc_hd__dlrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095000 0.415000 6.355000 2.455000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.500000 0.995000 5.435000 1.325000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 2.005000 ;
      RECT 2.715000  0.705000 3.095000 1.035000 ;
      RECT 2.840000  0.365000 3.500000 0.535000 ;
      RECT 2.900000  2.255000 3.650000 2.425000 ;
      RECT 2.925000  1.035000 3.095000 1.415000 ;
      RECT 2.925000  1.415000 3.265000 1.995000 ;
      RECT 3.330000  0.535000 3.500000 1.025000 ;
      RECT 3.330000  1.025000 4.330000 1.245000 ;
      RECT 3.480000  1.245000 4.330000 1.325000 ;
      RECT 3.480000  1.325000 3.650000 2.255000 ;
      RECT 3.740000  0.085000 4.070000 0.530000 ;
      RECT 3.820000  1.535000 5.925000 1.865000 ;
      RECT 3.820000  2.135000 4.110000 2.635000 ;
      RECT 4.240000  0.255000 4.590000 0.655000 ;
      RECT 4.240000  0.655000 5.925000 0.825000 ;
      RECT 4.300000  2.135000 4.580000 2.635000 ;
      RECT 4.750000  1.865000 4.940000 2.465000 ;
      RECT 5.095000  0.085000 5.925000 0.485000 ;
      RECT 5.110000  2.135000 5.925000 2.635000 ;
      RECT 5.605000  0.825000 5.925000 1.535000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.785000 2.640000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.445000 3.100000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.160000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.700000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 1.415000 3.160000 1.460000 ;
      RECT 2.870000 1.600000 3.160000 1.645000 ;
  END
END sky130_fd_sc_hd__dlrtn_1
MACRO sky130_fd_sc_hd__dlrtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.595000 0.255000 5.925000 0.485000 ;
        RECT 5.655000 1.875000 5.925000 2.465000 ;
        RECT 5.755000 0.485000 5.925000 0.765000 ;
        RECT 5.755000 0.765000 6.355000 0.865000 ;
        RECT 5.755000 1.425000 6.355000 1.500000 ;
        RECT 5.755000 1.500000 5.925000 1.875000 ;
        RECT 5.760000 1.415000 6.355000 1.425000 ;
        RECT 5.765000 1.410000 6.355000 1.415000 ;
        RECT 5.770000 0.865000 6.355000 0.890000 ;
        RECT 5.775000 1.385000 6.355000 1.410000 ;
        RECT 5.785000 0.890000 6.355000 1.385000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.480000 0.995000 5.170000 1.325000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.960000  0.785000 2.340000 1.095000 ;
      RECT 1.960000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 2.005000 ;
      RECT 2.675000  0.705000 3.095000 1.145000 ;
      RECT 2.775000  2.255000 3.605000 2.425000 ;
      RECT 2.810000  0.365000 3.500000 0.535000 ;
      RECT 2.925000  1.145000 3.095000 1.415000 ;
      RECT 2.925000  1.415000 3.265000 1.995000 ;
      RECT 3.330000  0.535000 3.500000 1.025000 ;
      RECT 3.330000  1.025000 4.310000 1.245000 ;
      RECT 3.435000  1.245000 4.310000 1.325000 ;
      RECT 3.435000  1.325000 3.605000 2.255000 ;
      RECT 3.735000  0.085000 4.070000 0.530000 ;
      RECT 3.800000  2.135000 4.110000 2.635000 ;
      RECT 3.820000  1.535000 5.585000 1.705000 ;
      RECT 3.820000  1.705000 4.920000 1.865000 ;
      RECT 4.240000  0.255000 4.590000 0.655000 ;
      RECT 4.240000  0.655000 5.585000 0.825000 ;
      RECT 4.280000  2.135000 4.560000 2.635000 ;
      RECT 4.730000  1.865000 4.920000 2.465000 ;
      RECT 5.090000  1.875000 5.460000 2.635000 ;
      RECT 5.095000  0.085000 5.425000 0.485000 ;
      RECT 5.350000  0.995000 5.615000 1.325000 ;
      RECT 5.415000  0.825000 5.585000 0.995000 ;
      RECT 5.415000  1.325000 5.585000 1.535000 ;
      RECT 6.095000  0.085000 6.355000 0.595000 ;
      RECT 6.095000  1.670000 6.355000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.785000 2.640000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.445000 3.100000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.160000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.700000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 1.415000 3.160000 1.460000 ;
      RECT 2.870000 1.600000 3.160000 1.645000 ;
  END
END sky130_fd_sc_hd__dlrtn_2
MACRO sky130_fd_sc_hd__dlrtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.955000 1.795000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.014750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.610000 0.255000 5.965000 0.485000 ;
        RECT 5.680000 1.875000 5.965000 2.465000 ;
        RECT 5.795000 0.485000 5.965000 0.765000 ;
        RECT 5.795000 0.765000 7.275000 1.325000 ;
        RECT 5.795000 1.325000 5.965000 1.875000 ;
        RECT 6.575000 0.255000 6.775000 0.765000 ;
        RECT 6.575000 1.325000 6.775000 2.465000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505000 0.995000 5.145000 1.325000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.360000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.960000 1.835000 2.275000 2.635000 ;
        RECT 3.825000 2.135000 4.115000 2.635000 ;
        RECT 4.305000 2.135000 4.585000 2.635000 ;
        RECT 5.115000 1.875000 5.485000 2.635000 ;
        RECT 6.135000 1.495000 6.405000 2.635000 ;
        RECT 6.945000 1.495000 7.275000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.460000  1.495000 2.145000 1.665000 ;
      RECT 1.460000  1.665000 1.790000 2.415000 ;
      RECT 1.540000  0.345000 1.710000 0.615000 ;
      RECT 1.540000  0.615000 2.145000 0.765000 ;
      RECT 1.540000  0.765000 2.345000 0.785000 ;
      RECT 1.880000  0.085000 2.210000 0.445000 ;
      RECT 1.975000  0.785000 2.345000 1.095000 ;
      RECT 1.975000  1.095000 2.145000 1.495000 ;
      RECT 2.475000  1.355000 2.760000 2.005000 ;
      RECT 2.720000  0.705000 3.100000 1.035000 ;
      RECT 2.845000  0.365000 3.505000 0.535000 ;
      RECT 2.905000  2.255000 3.655000 2.425000 ;
      RECT 2.930000  1.035000 3.100000 1.415000 ;
      RECT 2.930000  1.415000 3.270000 1.995000 ;
      RECT 3.335000  0.535000 3.505000 1.025000 ;
      RECT 3.335000  1.025000 4.315000 1.245000 ;
      RECT 3.485000  1.245000 4.315000 1.325000 ;
      RECT 3.485000  1.325000 3.655000 2.255000 ;
      RECT 3.745000  0.085000 4.075000 0.530000 ;
      RECT 3.825000  1.535000 5.625000 1.705000 ;
      RECT 3.825000  1.705000 4.945000 1.865000 ;
      RECT 4.245000  0.255000 4.595000 0.655000 ;
      RECT 4.245000  0.655000 5.625000 0.825000 ;
      RECT 4.755000  1.865000 4.945000 2.465000 ;
      RECT 5.100000  0.085000 5.440000 0.485000 ;
      RECT 5.455000  0.825000 5.625000 1.535000 ;
      RECT 6.135000  0.085000 6.405000 0.595000 ;
      RECT 6.945000  0.085000 7.275000 0.595000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.475000  1.785000 2.645000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.935000  1.445000 3.105000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.165000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.705000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.415000 1.755000 2.705000 1.800000 ;
      RECT 2.415000 1.940000 2.705000 1.985000 ;
      RECT 2.875000 1.415000 3.165000 1.460000 ;
      RECT 2.875000 1.600000 3.165000 1.645000 ;
  END
END sky130_fd_sc_hd__dlrtn_4
MACRO sky130_fd_sc_hd__dlrbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.536250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.650000 0.415000 5.910000 0.655000 ;
        RECT 5.650000 0.655000 5.950000 0.685000 ;
        RECT 5.650000 0.685000 5.975000 0.825000 ;
        RECT 5.650000 1.495000 5.975000 1.660000 ;
        RECT 5.650000 1.660000 5.915000 2.465000 ;
        RECT 5.740000 0.825000 5.975000 0.860000 ;
        RECT 5.790000 0.860000 5.975000 0.885000 ;
        RECT 5.790000 0.885000 6.355000 1.325000 ;
        RECT 5.790000 1.325000 5.975000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.500000 0.255000 7.755000 0.825000 ;
        RECT 7.500000 1.445000 7.755000 2.465000 ;
        RECT 7.545000 0.825000 7.755000 1.055000 ;
        RECT 7.545000 1.055000 8.195000 1.325000 ;
        RECT 7.545000 1.325000 7.755000 1.445000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.390000 0.995000 5.140000 1.325000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.780000 0.805000 ;
      RECT 0.085000  1.795000 0.780000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.605000  0.805000 0.780000 1.070000 ;
      RECT 0.605000  1.070000 0.840000 1.400000 ;
      RECT 0.605000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 2.005000 ;
      RECT 2.715000  0.705000 3.095000 1.035000 ;
      RECT 2.840000  0.365000 3.500000 0.535000 ;
      RECT 2.900000  2.255000 3.650000 2.425000 ;
      RECT 2.925000  1.035000 3.095000 1.415000 ;
      RECT 2.925000  1.415000 3.265000 1.995000 ;
      RECT 3.330000  0.535000 3.500000 0.995000 ;
      RECT 3.330000  0.995000 4.200000 1.165000 ;
      RECT 3.480000  1.165000 4.200000 1.325000 ;
      RECT 3.480000  1.325000 3.650000 2.255000 ;
      RECT 3.740000  0.085000 4.070000 0.825000 ;
      RECT 3.820000  2.135000 4.590000 2.635000 ;
      RECT 3.840000  1.495000 5.480000 1.665000 ;
      RECT 3.840000  1.665000 4.930000 1.865000 ;
      RECT 4.340000  0.415000 4.560000 0.655000 ;
      RECT 4.340000  0.655000 5.480000 0.825000 ;
      RECT 4.760000  1.865000 4.930000 2.435000 ;
      RECT 5.100000  0.085000 5.480000 0.485000 ;
      RECT 5.100000  1.855000 5.350000 2.635000 ;
      RECT 5.310000  0.825000 5.480000 0.995000 ;
      RECT 5.310000  0.995000 5.620000 1.325000 ;
      RECT 5.310000  1.325000 5.480000 1.495000 ;
      RECT 6.085000  0.085000 6.355000 0.545000 ;
      RECT 6.085000  1.830000 6.355000 2.635000 ;
      RECT 6.525000  0.255000 6.855000 0.995000 ;
      RECT 6.525000  0.995000 7.375000 1.325000 ;
      RECT 6.525000  1.325000 6.855000 2.465000 ;
      RECT 7.025000  0.085000 7.330000 0.545000 ;
      RECT 7.035000  1.835000 7.330000 2.635000 ;
      RECT 7.925000  0.085000 8.195000 0.885000 ;
      RECT 7.925000  1.495000 8.195000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.785000 2.640000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.445000 3.100000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.160000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.700000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 1.415000 3.160000 1.460000 ;
      RECT 2.870000 1.600000 3.160000 1.645000 ;
  END
END sky130_fd_sc_hd__dlrbn_2
MACRO sky130_fd_sc_hd__dlrbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.060000 0.255000 6.380000 2.465000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.475000 0.255000 7.735000 0.595000 ;
        RECT 7.475000 1.785000 7.735000 2.465000 ;
        RECT 7.560000 0.595000 7.735000 1.785000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.470000 0.995000 5.455000 1.325000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.780000 0.805000 ;
      RECT 0.085000  1.795000 0.780000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 2.005000 ;
      RECT 2.715000  0.705000 3.095000 1.035000 ;
      RECT 2.840000  0.365000 3.500000 0.535000 ;
      RECT 2.900000  2.255000 3.650000 2.425000 ;
      RECT 2.925000  1.035000 3.095000 1.415000 ;
      RECT 2.925000  1.415000 3.265000 1.995000 ;
      RECT 3.330000  0.535000 3.500000 0.995000 ;
      RECT 3.330000  0.995000 4.300000 1.165000 ;
      RECT 3.480000  1.165000 4.300000 1.325000 ;
      RECT 3.480000  1.325000 3.650000 2.255000 ;
      RECT 3.740000  0.085000 4.070000 0.530000 ;
      RECT 3.820000  2.135000 4.090000 2.635000 ;
      RECT 3.840000  1.535000 5.875000 1.765000 ;
      RECT 3.840000  1.765000 4.970000 1.865000 ;
      RECT 4.240000  0.255000 4.540000 0.655000 ;
      RECT 4.240000  0.655000 5.875000 0.825000 ;
      RECT 4.260000  2.135000 4.590000 2.635000 ;
      RECT 4.760000  1.865000 4.970000 2.435000 ;
      RECT 5.135000  0.085000 5.875000 0.485000 ;
      RECT 5.150000  1.935000 5.890000 2.635000 ;
      RECT 5.625000  0.825000 5.875000 1.535000 ;
      RECT 6.580000  0.255000 6.750000 0.985000 ;
      RECT 6.580000  0.985000 6.830000 0.995000 ;
      RECT 6.580000  0.995000 7.390000 1.325000 ;
      RECT 6.580000  1.325000 6.830000 2.465000 ;
      RECT 6.975000  0.085000 7.305000 0.465000 ;
      RECT 7.010000  1.835000 7.305000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.785000 2.640000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.445000 3.100000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.160000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.700000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 1.415000 3.160000 1.460000 ;
      RECT 2.870000 1.600000 3.160000 1.645000 ;
  END
END sky130_fd_sc_hd__dlrbn_1
MACRO sky130_fd_sc_hd__o22a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095000 1.075000 3.590000 1.275000 ;
        RECT 3.270000 1.275000 3.590000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.595000 1.075000 2.925000 1.325000 ;
        RECT 2.745000 1.325000 2.925000 1.445000 ;
        RECT 2.745000 1.445000 3.100000 1.615000 ;
        RECT 2.900000 1.615000 3.100000 2.405000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 1.075000 1.790000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 1.075000 2.425000 1.325000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 0.365000 0.805000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.130000 -0.085000 0.300000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.115000  1.445000 0.365000 2.635000 ;
      RECT 0.185000  0.085000 0.355000 0.885000 ;
      RECT 0.975000  0.715000 2.215000 0.895000 ;
      RECT 0.975000  0.895000 1.255000 1.495000 ;
      RECT 0.975000  1.495000 2.575000 1.705000 ;
      RECT 0.995000  1.875000 1.795000 2.635000 ;
      RECT 1.025000  0.085000 1.205000 0.545000 ;
      RECT 1.465000  0.295000 2.730000 0.475000 ;
      RECT 1.850000  0.645000 2.215000 0.715000 ;
      RECT 2.190000  1.705000 2.575000 2.465000 ;
      RECT 2.390000  0.475000 2.730000 0.695000 ;
      RECT 2.390000  0.695000 3.590000 0.825000 ;
      RECT 2.560000  0.825000 3.590000 0.865000 ;
      RECT 2.915000  0.085000 3.085000 0.525000 ;
      RECT 3.255000  0.280000 3.590000 0.695000 ;
      RECT 3.270000  1.795000 3.590000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o22a_2
MACRO sky130_fd_sc_hd__o22a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.670000 1.075000 3.135000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.165000 1.075000 2.495000 1.325000 ;
        RECT 2.315000 1.325000 2.495000 1.445000 ;
        RECT 2.315000 1.445000 2.645000 1.615000 ;
        RECT 2.445000 1.615000 2.645000 2.405000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.980000 1.075000 1.335000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 1.075000 1.995000 1.325000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.365000 0.365000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.535000  0.715000 1.785000 0.895000 ;
      RECT 0.535000  0.895000 0.810000 1.495000 ;
      RECT 0.535000  1.495000 2.145000 1.705000 ;
      RECT 0.555000  1.875000 1.340000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 1.035000  0.295000 2.285000 0.475000 ;
      RECT 1.420000  0.645000 1.785000 0.715000 ;
      RECT 1.735000  1.705000 2.145000 1.805000 ;
      RECT 1.735000  1.805000 2.120000 2.465000 ;
      RECT 1.955000  0.475000 2.285000 0.695000 ;
      RECT 1.955000  0.695000 3.135000 0.865000 ;
      RECT 2.455000  0.085000 2.625000 0.525000 ;
      RECT 2.795000  0.280000 3.135000 0.695000 ;
      RECT 2.815000  1.455000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o22a_1
MACRO sky130_fd_sc_hd__o22a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.350000 1.075000 4.680000 1.445000 ;
        RECT 4.350000 1.445000 5.735000 1.615000 ;
        RECT 5.565000 1.075000 6.355000 1.275000 ;
        RECT 5.565000 1.275000 5.735000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.900000 1.075000 5.395000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.420000 1.075000 2.955000 1.445000 ;
        RECT 2.420000 1.445000 4.180000 1.615000 ;
        RECT 3.850000 1.075000 4.180000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.125000 1.075000 3.680000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.725000 1.770000 0.905000 ;
        RECT 0.085000 0.905000 0.370000 1.445000 ;
        RECT 0.085000 1.445000 1.730000 1.615000 ;
        RECT 0.600000 0.265000 0.930000 0.725000 ;
        RECT 0.640000 1.615000 0.890000 2.465000 ;
        RECT 1.440000 0.255000 1.770000 0.725000 ;
        RECT 1.480000 1.615000 1.730000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.220000  1.825000 0.470000 2.635000 ;
      RECT 0.260000  0.085000 0.430000 0.555000 ;
      RECT 0.540000  1.075000 2.230000 1.275000 ;
      RECT 1.060000  1.795000 1.310000 2.635000 ;
      RECT 1.100000  0.085000 1.270000 0.555000 ;
      RECT 1.900000  1.275000 2.230000 1.785000 ;
      RECT 1.900000  1.785000 5.270000 1.955000 ;
      RECT 1.900000  2.125000 2.670000 2.635000 ;
      RECT 1.940000  0.085000 2.110000 0.555000 ;
      RECT 1.940000  0.735000 3.970000 0.905000 ;
      RECT 1.940000  0.905000 2.230000 1.075000 ;
      RECT 2.380000  0.255000 4.470000 0.475000 ;
      RECT 2.415000  0.645000 3.970000 0.735000 ;
      RECT 2.840000  2.125000 3.090000 2.295000 ;
      RECT 2.840000  2.295000 3.930000 2.465000 ;
      RECT 3.260000  1.955000 3.510000 2.125000 ;
      RECT 3.680000  2.125000 3.930000 2.295000 ;
      RECT 4.100000  2.125000 4.430000 2.635000 ;
      RECT 4.140000  0.475000 4.470000 0.735000 ;
      RECT 4.140000  0.735000 6.150000 0.905000 ;
      RECT 4.600000  2.125000 4.850000 2.295000 ;
      RECT 4.600000  2.295000 5.690000 2.465000 ;
      RECT 4.640000  0.085000 4.810000 0.555000 ;
      RECT 4.980000  0.255000 5.310000 0.725000 ;
      RECT 4.980000  0.725000 6.150000 0.735000 ;
      RECT 5.020000  1.955000 5.270000 2.125000 ;
      RECT 5.440000  1.785000 5.690000 2.295000 ;
      RECT 5.480000  0.085000 5.650000 0.555000 ;
      RECT 5.820000  0.255000 6.150000 0.725000 ;
      RECT 5.905000  1.455000 6.110000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__o22a_4
MACRO sky130_fd_sc_hd__probec_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__probec_p_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.240000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT -1.140000 0.770000 0.040000 1.950000 ;
        RECT  1.460000 0.770000 2.640000 1.950000 ;
    END
    PORT
      LAYER met5 ;
        RECT -1.260000  0.560000 2.760000 2.160000 ;
        RECT  1.160000 -1.105000 2.760000 0.560000 ;
        RECT  1.160000  2.160000 2.760000 3.825000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 4.360000 -1.170000 6.675000 0.560000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 4.360000 2.160000 6.675000 3.890000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.095000  1.445000 1.595000 1.615000 ;
      RECT 0.095000  1.615000 0.425000 2.465000 ;
      RECT 0.175000  0.255000 0.345000 0.735000 ;
      RECT 0.175000  0.735000 1.595000 0.905000 ;
      RECT 0.515000  0.085000 0.845000 0.565000 ;
      RECT 0.595000  1.835000 0.765000 2.635000 ;
      RECT 0.935000  1.615000 1.265000 2.465000 ;
      RECT 1.015000  0.260000 1.185000 0.735000 ;
      RECT 1.355000  0.085000 1.685000 0.565000 ;
      RECT 1.420000  0.905000 1.595000 1.075000 ;
      RECT 1.420000  1.075000 4.045000 1.245000 ;
      RECT 1.420000  1.245000 1.595000 1.445000 ;
      RECT 1.435000  1.835000 1.605000 2.635000 ;
      RECT 1.855000  0.255000 2.025000 0.735000 ;
      RECT 1.855000  0.735000 4.545000 0.905000 ;
      RECT 1.855000  1.445000 4.545000 1.615000 ;
      RECT 1.855000  1.615000 2.025000 2.465000 ;
      RECT 2.195000  0.085000 2.525000 0.565000 ;
      RECT 2.195000  1.835000 2.525000 2.635000 ;
      RECT 2.695000  0.255000 2.865000 0.735000 ;
      RECT 2.695000  1.615000 2.865000 2.465000 ;
      RECT 3.035000  0.085000 3.365000 0.565000 ;
      RECT 3.035000  1.835000 3.365000 2.635000 ;
      RECT 3.535000  0.255000 3.705000 0.735000 ;
      RECT 3.535000  1.615000 3.705000 2.465000 ;
      RECT 3.875000  0.085000 4.205000 0.565000 ;
      RECT 3.875000  1.835000 4.205000 2.635000 ;
      RECT 4.290000  0.905000 4.545000 1.055000 ;
      RECT 4.290000  1.055000 4.870000 1.315000 ;
      RECT 4.290000  1.315000 4.545000 1.445000 ;
      RECT 4.375000  0.255000 4.545000 0.735000 ;
      RECT 4.375000  1.615000 4.545000 2.465000 ;
      RECT 4.715000  0.085000 5.045000 0.885000 ;
      RECT 4.715000  1.485000 5.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.305000  1.105000 4.475000 1.275000 ;
      RECT 4.665000  1.105000 4.835000 1.275000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 5.520000 -0.130000 ;
      RECT 0.000000 -0.130000 5.840000  0.130000 ;
      RECT 0.000000  0.130000 5.520000  0.240000 ;
      RECT 0.000000  2.480000 5.520000  2.590000 ;
      RECT 0.000000  2.590000 5.840000  2.850000 ;
      RECT 0.000000  2.850000 5.520000  2.960000 ;
      RECT 2.020000  1.060000 2.660000  1.120000 ;
      RECT 2.020000  1.120000 4.895000  1.260000 ;
      RECT 2.020000  1.260000 2.660000  1.320000 ;
      RECT 4.245000  1.075000 4.895000  1.120000 ;
      RECT 4.245000  1.260000 4.895000  1.305000 ;
    LAYER met2 ;
      RECT 1.890000  1.050000 2.660000 1.330000 ;
      RECT 5.135000 -0.140000 5.905000 0.140000 ;
      RECT 5.135000  2.580000 5.905000 2.860000 ;
    LAYER met3 ;
      RECT -0.715000  1.030000 0.065000 1.350000 ;
      RECT  1.885000  1.025000 2.665000 1.355000 ;
      RECT  5.130000 -0.165000 5.910000 0.165000 ;
      RECT  5.130000  2.555000 5.910000 2.885000 ;
    LAYER met4 ;
      RECT 4.930000 -0.895000 6.110000 0.285000 ;
      RECT 4.930000  2.435000 6.110000 3.615000 ;
    LAYER via ;
      RECT 2.050000  1.060000 2.310000 1.320000 ;
      RECT 2.370000  1.060000 2.630000 1.320000 ;
      RECT 5.230000 -0.130000 5.490000 0.130000 ;
      RECT 5.230000  2.590000 5.490000 2.850000 ;
      RECT 5.550000 -0.130000 5.810000 0.130000 ;
      RECT 5.550000  2.590000 5.810000 2.850000 ;
    LAYER via2 ;
      RECT 1.935000  1.050000 2.215000 1.330000 ;
      RECT 2.335000  1.050000 2.615000 1.330000 ;
      RECT 5.180000 -0.140000 5.460000 0.140000 ;
      RECT 5.180000  2.580000 5.460000 2.860000 ;
      RECT 5.580000 -0.140000 5.860000 0.140000 ;
      RECT 5.580000  2.580000 5.860000 2.860000 ;
    LAYER via3 ;
      RECT -0.685000  1.030000 -0.365000 1.350000 ;
      RECT -0.285000  1.030000  0.035000 1.350000 ;
      RECT  1.915000  1.030000  2.235000 1.350000 ;
      RECT  2.315000  1.030000  2.635000 1.350000 ;
      RECT  5.160000 -0.160000  5.480000 0.160000 ;
      RECT  5.160000  2.560000  5.480000 2.880000 ;
      RECT  5.560000 -0.160000  5.880000 0.160000 ;
      RECT  5.560000  2.560000  5.880000 2.880000 ;
  END
END sky130_fd_sc_hd__probec_p_8
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.072500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.255000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 1.085000 ;
        RECT 5.360000 1.085000 6.555000 1.410000 ;
        RECT 5.360000 1.410000 5.635000 2.370000 ;
        RECT 6.280000 1.410000 6.555000 2.370000 ;
        RECT 6.335000 0.255000 6.555000 1.085000 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 7.290000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 7.360000 5.680000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.075000 5.245000 0.200000 5.395000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.250000 1.305000 7.405000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 7.360000 5.525000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.255000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.255000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 7.360000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.825000  0.085000 6.155000 0.845000 ;
      RECT 5.905000  1.610000 6.075000 2.635000 ;
      RECT 6.755000  0.085000 7.005000 0.925000 ;
      RECT 6.755000  1.610000 6.935000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.585000  5.355000 6.755000 5.525000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.045000  5.355000 7.215000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 7.360000 0.240000 ;
    LAYER nwell ;
      RECT -0.190000 1.305000 0.650000 4.135000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4
MACRO sky130_fd_sc_hd__sedfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.80000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755000 0.305000 13.085000 2.420000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 1.105000 6.215000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.105000 5.250000 1.615000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.800000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  4.885000 1.435000 ;
        RECT -0.190000 1.435000 13.990000 2.910000 ;
        RECT  7.200000 1.305000 13.990000 1.435000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.800000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.800000 0.085000 ;
      RECT  0.000000  2.635000 13.800000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.595000  0.255000  4.795000 0.645000 ;
      RECT  4.595000  0.645000  4.855000 0.825000 ;
      RECT  4.635000  2.210000  4.965000 2.465000 ;
      RECT  4.685000  0.825000  4.855000 1.785000 ;
      RECT  4.685000  1.785000  4.965000 2.210000 ;
      RECT  4.965000  0.255000  5.590000 0.515000 ;
      RECT  5.155000  1.835000  6.585000 2.005000 ;
      RECT  5.155000  2.005000  5.495000 2.465000 ;
      RECT  5.260000  0.515000  5.590000 0.935000 ;
      RECT  5.420000  0.935000  5.590000 1.835000 ;
      RECT  5.665000  2.175000  6.010000 2.635000 ;
      RECT  5.760000  0.085000  6.010000 0.905000 ;
      RECT  6.385000  1.355000  6.585000 1.835000 ;
      RECT  6.515000  0.255000  7.135000 0.565000 ;
      RECT  6.515000  0.565000  6.925000 1.185000 ;
      RECT  6.675000  2.150000  7.005000 2.465000 ;
      RECT  6.755000  1.185000  6.925000 1.865000 ;
      RECT  6.755000  1.865000  7.005000 2.150000 ;
      RECT  7.095000  1.125000  7.280000 1.720000 ;
      RECT  7.115000  0.735000  7.620000 0.955000 ;
      RECT  7.215000  2.175000  8.255000 2.375000 ;
      RECT  7.305000  0.255000  7.980000 0.565000 ;
      RECT  7.450000  0.955000  7.620000 1.655000 ;
      RECT  7.450000  1.655000  7.915000 2.005000 ;
      RECT  7.810000  0.565000  7.980000 1.315000 ;
      RECT  7.810000  1.315000  8.660000 1.485000 ;
      RECT  8.085000  1.485000  8.660000 1.575000 ;
      RECT  8.085000  1.575000  8.255000 2.175000 ;
      RECT  8.170000  0.765000  9.235000 1.045000 ;
      RECT  8.170000  1.045000  9.745000 1.065000 ;
      RECT  8.170000  1.065000  8.370000 1.095000 ;
      RECT  8.245000  0.085000  8.640000 0.560000 ;
      RECT  8.425000  1.835000  8.660000 2.635000 ;
      RECT  8.490000  1.245000  8.660000 1.315000 ;
      RECT  8.830000  0.255000  9.235000 0.765000 ;
      RECT  8.830000  1.065000  9.745000 1.375000 ;
      RECT  8.830000  1.375000  9.160000 2.465000 ;
      RECT  9.370000  2.105000  9.660000 2.635000 ;
      RECT  9.465000  0.085000  9.740000 0.615000 ;
      RECT 10.090000  1.245000 10.280000 1.965000 ;
      RECT 10.225000  2.165000 11.110000 2.355000 ;
      RECT 10.305000  0.705000 10.770000 1.035000 ;
      RECT 10.325000  0.330000 11.110000 0.535000 ;
      RECT 10.450000  1.035000 10.770000 1.995000 ;
      RECT 10.940000  0.535000 11.110000 0.995000 ;
      RECT 10.940000  0.995000 11.810000 1.325000 ;
      RECT 10.940000  1.325000 11.110000 2.165000 ;
      RECT 11.280000  1.530000 12.180000 1.905000 ;
      RECT 11.280000  2.135000 11.540000 2.635000 ;
      RECT 11.350000  0.085000 11.665000 0.615000 ;
      RECT 11.840000  1.905000 12.180000 2.465000 ;
      RECT 11.850000  0.300000 12.180000 0.825000 ;
      RECT 11.990000  0.825000 12.180000 1.530000 ;
      RECT 12.350000  0.085000 12.585000 0.900000 ;
      RECT 12.350000  1.465000 12.585000 2.635000 ;
      RECT 13.255000  0.085000 13.515000 0.900000 ;
      RECT 13.255000  1.465000 13.515000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.615000  0.425000  4.785000 0.595000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.530000  0.425000  6.700000 0.595000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.100000  1.445000  7.270000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.510000  1.785000  7.680000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.100000  1.785000 10.270000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.520000  1.445000 10.690000 1.615000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.000000  0.765000 12.170000 0.935000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000 10.330000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000 10.750000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 12.230000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.555000 0.395000  6.760000 0.580000 ;
      RECT  4.555000 0.580000  4.845000 0.625000 ;
      RECT  6.470000 0.580000  6.760000 0.625000 ;
      RECT  7.040000 1.415000  7.330000 1.460000 ;
      RECT  7.040000 1.600000  7.330000 1.645000 ;
      RECT  7.450000 1.755000  7.740000 1.800000 ;
      RECT  7.450000 1.940000  7.740000 1.985000 ;
      RECT 10.040000 1.755000 10.330000 1.800000 ;
      RECT 10.040000 1.940000 10.330000 1.985000 ;
      RECT 10.460000 1.415000 10.750000 1.460000 ;
      RECT 10.460000 1.600000 10.750000 1.645000 ;
      RECT 11.940000 0.735000 12.230000 0.780000 ;
      RECT 11.940000 0.920000 12.230000 0.965000 ;
  END
END sky130_fd_sc_hd__sedfxtp_2
MACRO sky130_fd_sc_hd__sedfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.72000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755000 0.305000 13.085000 1.070000 ;
        RECT 12.755000 1.070000 13.925000 1.295000 ;
        RECT 12.755000 1.295000 13.085000 2.420000 ;
        RECT 13.595000 0.305000 13.925000 1.070000 ;
        RECT 13.595000 1.295000 13.925000 2.420000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 1.105000 6.215000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.105000 5.250000 1.615000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.720000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  4.885000 1.435000 ;
        RECT -0.190000 1.435000 14.910000 2.910000 ;
        RECT  7.200000 1.305000 14.910000 1.435000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.720000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.720000 0.085000 ;
      RECT  0.000000  2.635000 14.720000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.595000  0.255000  4.795000 0.645000 ;
      RECT  4.595000  0.645000  4.855000 0.825000 ;
      RECT  4.635000  2.210000  4.965000 2.465000 ;
      RECT  4.685000  0.825000  4.855000 1.785000 ;
      RECT  4.685000  1.785000  4.965000 2.210000 ;
      RECT  4.965000  0.255000  5.590000 0.515000 ;
      RECT  5.155000  1.835000  6.585000 2.005000 ;
      RECT  5.155000  2.005000  5.495000 2.465000 ;
      RECT  5.260000  0.515000  5.590000 0.935000 ;
      RECT  5.420000  0.935000  5.590000 1.835000 ;
      RECT  5.665000  2.175000  6.010000 2.635000 ;
      RECT  5.760000  0.085000  6.010000 0.905000 ;
      RECT  6.385000  1.355000  6.585000 1.835000 ;
      RECT  6.515000  0.255000  7.135000 0.565000 ;
      RECT  6.515000  0.565000  6.925000 1.185000 ;
      RECT  6.675000  2.150000  7.005000 2.465000 ;
      RECT  6.755000  1.185000  6.925000 1.865000 ;
      RECT  6.755000  1.865000  7.005000 2.150000 ;
      RECT  7.095000  1.125000  7.280000 1.720000 ;
      RECT  7.115000  0.735000  7.620000 0.955000 ;
      RECT  7.215000  2.175000  8.255000 2.375000 ;
      RECT  7.305000  0.255000  7.980000 0.565000 ;
      RECT  7.450000  0.955000  7.620000 1.655000 ;
      RECT  7.450000  1.655000  7.915000 2.005000 ;
      RECT  7.810000  0.565000  7.980000 1.315000 ;
      RECT  7.810000  1.315000  8.660000 1.485000 ;
      RECT  8.085000  1.485000  8.660000 1.575000 ;
      RECT  8.085000  1.575000  8.255000 2.175000 ;
      RECT  8.170000  0.765000  9.235000 1.045000 ;
      RECT  8.170000  1.045000  9.745000 1.065000 ;
      RECT  8.170000  1.065000  8.370000 1.095000 ;
      RECT  8.245000  0.085000  8.640000 0.560000 ;
      RECT  8.425000  1.835000  8.660000 2.635000 ;
      RECT  8.490000  1.245000  8.660000 1.315000 ;
      RECT  8.830000  0.255000  9.235000 0.765000 ;
      RECT  8.830000  1.065000  9.745000 1.375000 ;
      RECT  8.830000  1.375000  9.160000 2.465000 ;
      RECT  9.370000  2.105000  9.660000 2.635000 ;
      RECT  9.465000  0.085000  9.740000 0.615000 ;
      RECT 10.090000  1.245000 10.280000 1.965000 ;
      RECT 10.225000  2.165000 11.110000 2.355000 ;
      RECT 10.305000  0.705000 10.770000 1.035000 ;
      RECT 10.325000  0.330000 11.110000 0.535000 ;
      RECT 10.450000  1.035000 10.770000 1.995000 ;
      RECT 10.940000  0.535000 11.110000 0.995000 ;
      RECT 10.940000  0.995000 11.810000 1.325000 ;
      RECT 10.940000  1.325000 11.110000 2.165000 ;
      RECT 11.280000  1.530000 12.180000 1.905000 ;
      RECT 11.280000  2.135000 11.540000 2.635000 ;
      RECT 11.350000  0.085000 11.665000 0.615000 ;
      RECT 11.840000  1.905000 12.180000 2.465000 ;
      RECT 11.850000  0.300000 12.180000 0.825000 ;
      RECT 11.990000  0.825000 12.180000 1.530000 ;
      RECT 12.350000  0.085000 12.585000 0.900000 ;
      RECT 12.350000  1.465000 12.585000 2.635000 ;
      RECT 13.255000  0.085000 13.425000 0.900000 ;
      RECT 13.255000  1.465000 13.425000 2.635000 ;
      RECT 14.095000  0.085000 14.355000 1.280000 ;
      RECT 14.095000  1.465000 14.355000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.615000  0.425000  4.785000 0.595000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.530000  0.425000  6.700000 0.595000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.100000  1.445000  7.270000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.510000  1.785000  7.680000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.100000  1.785000 10.270000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.520000  1.445000 10.690000 1.615000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.000000  0.765000 12.170000 0.935000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000 10.330000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000 10.750000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 12.230000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.555000 0.395000  6.760000 0.580000 ;
      RECT  4.555000 0.580000  4.845000 0.625000 ;
      RECT  6.470000 0.580000  6.760000 0.625000 ;
      RECT  7.040000 1.415000  7.330000 1.460000 ;
      RECT  7.040000 1.600000  7.330000 1.645000 ;
      RECT  7.450000 1.755000  7.740000 1.800000 ;
      RECT  7.450000 1.940000  7.740000 1.985000 ;
      RECT 10.040000 1.755000 10.330000 1.800000 ;
      RECT 10.040000 1.940000 10.330000 1.985000 ;
      RECT 10.460000 1.415000 10.750000 1.460000 ;
      RECT 10.460000 1.600000 10.750000 1.645000 ;
      RECT 11.940000 0.735000 12.230000 0.780000 ;
      RECT 11.940000 0.920000 12.230000 0.965000 ;
  END
END sky130_fd_sc_hd__sedfxtp_4
MACRO sky130_fd_sc_hd__sedfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.34000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.765000 0.305000 13.095000 2.420000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 1.105000 6.215000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.105000 5.250000 1.615000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  4.885000 1.435000 ;
        RECT -0.190000 1.435000 13.530000 2.910000 ;
        RECT  7.200000 1.305000 13.530000 1.435000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.340000 0.085000 ;
      RECT  0.000000  2.635000 13.340000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.595000  0.255000  4.795000 0.645000 ;
      RECT  4.595000  0.645000  4.855000 0.825000 ;
      RECT  4.635000  2.210000  4.965000 2.465000 ;
      RECT  4.685000  0.825000  4.855000 1.785000 ;
      RECT  4.685000  1.785000  4.965000 2.210000 ;
      RECT  4.965000  0.255000  5.590000 0.515000 ;
      RECT  5.155000  1.835000  6.585000 2.005000 ;
      RECT  5.155000  2.005000  5.495000 2.465000 ;
      RECT  5.260000  0.515000  5.590000 0.935000 ;
      RECT  5.420000  0.935000  5.590000 1.835000 ;
      RECT  5.665000  2.175000  6.010000 2.635000 ;
      RECT  5.760000  0.085000  6.010000 0.905000 ;
      RECT  6.385000  1.355000  6.585000 1.835000 ;
      RECT  6.515000  0.255000  7.135000 0.565000 ;
      RECT  6.515000  0.565000  6.925000 1.185000 ;
      RECT  6.675000  2.150000  7.005000 2.465000 ;
      RECT  6.755000  1.185000  6.925000 1.865000 ;
      RECT  6.755000  1.865000  7.005000 2.150000 ;
      RECT  7.095000  1.125000  7.280000 1.720000 ;
      RECT  7.115000  0.735000  7.620000 0.955000 ;
      RECT  7.215000  2.175000  8.255000 2.375000 ;
      RECT  7.305000  0.255000  7.980000 0.565000 ;
      RECT  7.450000  0.955000  7.620000 1.655000 ;
      RECT  7.450000  1.655000  7.915000 2.005000 ;
      RECT  7.810000  0.565000  7.980000 1.315000 ;
      RECT  7.810000  1.315000  8.660000 1.485000 ;
      RECT  8.085000  1.485000  8.660000 1.575000 ;
      RECT  8.085000  1.575000  8.255000 2.175000 ;
      RECT  8.170000  0.765000  9.235000 1.045000 ;
      RECT  8.170000  1.045000  9.745000 1.065000 ;
      RECT  8.170000  1.065000  8.370000 1.095000 ;
      RECT  8.245000  0.085000  8.640000 0.560000 ;
      RECT  8.425000  1.835000  8.660000 2.635000 ;
      RECT  8.490000  1.245000  8.660000 1.315000 ;
      RECT  8.830000  0.255000  9.235000 0.765000 ;
      RECT  8.830000  1.065000  9.745000 1.375000 ;
      RECT  8.830000  1.375000  9.160000 2.465000 ;
      RECT  9.370000  2.105000  9.660000 2.635000 ;
      RECT  9.465000  0.085000  9.740000 0.615000 ;
      RECT 10.090000  1.245000 10.280000 1.965000 ;
      RECT 10.225000  2.165000 11.110000 2.355000 ;
      RECT 10.305000  0.705000 10.770000 1.035000 ;
      RECT 10.325000  0.330000 11.110000 0.535000 ;
      RECT 10.450000  1.035000 10.770000 1.995000 ;
      RECT 10.940000  0.535000 11.110000 0.995000 ;
      RECT 10.940000  0.995000 11.810000 1.325000 ;
      RECT 10.940000  1.325000 11.110000 2.165000 ;
      RECT 11.280000  1.530000 12.180000 1.905000 ;
      RECT 11.280000  2.135000 11.540000 2.635000 ;
      RECT 11.350000  0.085000 11.665000 0.615000 ;
      RECT 11.840000  1.905000 12.180000 2.465000 ;
      RECT 11.850000  0.300000 12.180000 0.825000 ;
      RECT 11.990000  0.825000 12.180000 1.530000 ;
      RECT 12.350000  0.085000 12.595000 0.900000 ;
      RECT 12.350000  1.465000 12.595000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.615000  0.425000  4.785000 0.595000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.530000  0.425000  6.700000 0.595000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.100000  1.445000  7.270000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.510000  1.785000  7.680000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.100000  1.785000 10.270000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.520000  1.445000 10.690000 1.615000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.000000  0.765000 12.170000 0.935000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000 10.330000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000 10.750000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 12.230000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.555000 0.395000  6.760000 0.580000 ;
      RECT  4.555000 0.580000  4.845000 0.625000 ;
      RECT  6.470000 0.580000  6.760000 0.625000 ;
      RECT  7.040000 1.415000  7.330000 1.460000 ;
      RECT  7.040000 1.600000  7.330000 1.645000 ;
      RECT  7.450000 1.755000  7.740000 1.800000 ;
      RECT  7.450000 1.940000  7.740000 1.985000 ;
      RECT 10.040000 1.755000 10.330000 1.800000 ;
      RECT 10.040000 1.940000 10.330000 1.985000 ;
      RECT 10.460000 1.415000 10.750000 1.460000 ;
      RECT 10.460000 1.600000 10.750000 1.645000 ;
      RECT 11.940000 0.735000 12.230000 0.780000 ;
      RECT 11.940000 0.920000 12.230000 0.965000 ;
  END
END sky130_fd_sc_hd__sedfxtp_1
MACRO sky130_fd_sc_hd__dfbbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfbbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.88000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.760000 1.005000 2.170000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.115000 0.255000 12.345000 0.825000 ;
        RECT 12.115000 1.445000 12.345000 2.465000 ;
        RECT 12.160000 0.825000 12.345000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.240000 0.255000 10.500000 0.715000 ;
        RECT 10.240000 1.630000 10.500000 2.465000 ;
        RECT 10.320000 0.715000 10.500000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.250000 1.095000 9.730000 1.325000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.600000 0.735000 4.010000 0.965000 ;
        RECT 3.600000 0.965000 3.930000 1.065000 ;
      LAYER mcon ;
        RECT 3.840000 0.765000 4.010000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.470000 0.735000 7.845000 1.065000 ;
      LAYER mcon ;
        RECT 7.520000 0.765000 7.690000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.780000 0.735000 4.070000 0.780000 ;
        RECT 3.780000 0.780000 7.750000 0.920000 ;
        RECT 3.780000 0.920000 4.070000 0.965000 ;
        RECT 7.460000 0.735000 7.750000 0.780000 ;
        RECT 7.460000 0.920000 7.750000 0.965000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.440000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 13.070000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.880000 0.085000 ;
      RECT  0.000000  2.635000 12.880000 2.805000 ;
      RECT  0.085000  0.345000  0.345000 0.635000 ;
      RECT  0.085000  0.635000  0.840000 0.805000 ;
      RECT  0.085000  1.795000  0.840000 1.965000 ;
      RECT  0.085000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.240000 2.465000 ;
      RECT  1.420000  0.635000  2.125000 0.825000 ;
      RECT  1.420000  0.825000  1.590000 1.795000 ;
      RECT  1.420000  1.795000  2.125000 1.965000 ;
      RECT  1.445000  0.085000  1.785000 0.465000 ;
      RECT  1.445000  2.135000  1.785000 2.635000 ;
      RECT  1.955000  0.305000  2.125000 0.635000 ;
      RECT  1.955000  1.965000  2.125000 2.465000 ;
      RECT  2.340000  0.705000  2.560000 1.575000 ;
      RECT  2.340000  1.575000  2.840000 1.955000 ;
      RECT  2.350000  2.250000  3.180000 2.420000 ;
      RECT  2.415000  0.265000  3.410000 0.465000 ;
      RECT  2.740000  0.645000  3.070000 1.015000 ;
      RECT  3.010000  1.195000  3.410000 1.235000 ;
      RECT  3.010000  1.235000  4.360000 1.405000 ;
      RECT  3.010000  1.405000  3.180000 2.250000 ;
      RECT  3.240000  0.465000  3.410000 1.195000 ;
      RECT  3.350000  1.575000  3.600000 1.785000 ;
      RECT  3.350000  1.785000  4.700000 2.035000 ;
      RECT  3.420000  2.205000  3.800000 2.635000 ;
      RECT  3.580000  0.085000  3.750000 0.525000 ;
      RECT  3.920000  0.255000  5.170000 0.425000 ;
      RECT  3.920000  0.425000  4.250000 0.545000 ;
      RECT  4.100000  2.035000  4.270000 2.375000 ;
      RECT  4.110000  1.405000  4.360000 1.485000 ;
      RECT  4.140000  1.155000  4.360000 1.235000 ;
      RECT  4.420000  0.595000  4.750000 0.765000 ;
      RECT  4.530000  0.765000  4.750000 0.895000 ;
      RECT  4.530000  0.895000  5.840000 1.065000 ;
      RECT  4.530000  1.065000  4.700000 1.785000 ;
      RECT  4.870000  1.235000  5.200000 1.415000 ;
      RECT  4.870000  1.415000  5.875000 1.655000 ;
      RECT  4.890000  1.915000  5.220000 2.635000 ;
      RECT  4.920000  0.425000  5.170000 0.715000 ;
      RECT  5.360000  0.085000  5.690000 0.465000 ;
      RECT  5.510000  1.065000  5.840000 1.235000 ;
      RECT  6.075000  1.575000  6.310000 1.985000 ;
      RECT  6.135000  0.705000  6.420000 1.125000 ;
      RECT  6.135000  1.125000  6.755000 1.305000 ;
      RECT  6.265000  2.250000  7.095000 2.420000 ;
      RECT  6.330000  0.265000  7.095000 0.465000 ;
      RECT  6.550000  1.305000  6.755000 1.905000 ;
      RECT  6.925000  0.465000  7.095000 1.235000 ;
      RECT  6.925000  1.235000  8.275000 1.405000 ;
      RECT  6.925000  1.405000  7.095000 2.250000 ;
      RECT  7.265000  1.575000  7.515000 1.915000 ;
      RECT  7.265000  1.915000 10.070000 2.085000 ;
      RECT  7.275000  0.085000  7.535000 0.525000 ;
      RECT  7.335000  2.255000  7.715000 2.635000 ;
      RECT  7.795000  0.255000  8.965000 0.425000 ;
      RECT  7.795000  0.425000  8.125000 0.545000 ;
      RECT  7.955000  2.085000  8.125000 2.375000 ;
      RECT  8.055000  1.075000  8.275000 1.235000 ;
      RECT  8.295000  0.595000  8.625000 0.780000 ;
      RECT  8.445000  0.780000  8.625000 1.915000 ;
      RECT  8.655000  2.255000 10.070000 2.635000 ;
      RECT  8.795000  0.425000  8.965000 0.585000 ;
      RECT  8.795000  0.755000  9.500000 0.925000 ;
      RECT  8.795000  0.925000  9.070000 1.575000 ;
      RECT  8.795000  1.575000  9.570000 1.745000 ;
      RECT  9.280000  0.265000  9.500000 0.755000 ;
      RECT  9.740000  0.085000 10.070000 0.805000 ;
      RECT  9.900000  0.995000 10.140000 1.325000 ;
      RECT  9.900000  1.325000 10.070000 1.915000 ;
      RECT 10.680000  0.085000 10.910000 0.885000 ;
      RECT 10.680000  1.465000 10.910000 2.635000 ;
      RECT 11.215000  0.255000 11.470000 0.995000 ;
      RECT 11.215000  0.995000 11.990000 1.325000 ;
      RECT 11.215000  1.325000 11.470000 2.415000 ;
      RECT 11.650000  0.085000 11.945000 0.545000 ;
      RECT 11.650000  1.765000 11.945000 2.635000 ;
      RECT 12.515000  0.085000 12.795000 0.885000 ;
      RECT 12.515000  1.465000 12.795000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.610000  0.765000  0.780000 0.935000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.070000  1.785000  1.240000 1.955000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.460000  1.785000  2.630000 1.955000 ;
      RECT  2.900000  0.765000  3.070000 0.935000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.680000  1.445000  5.850000 1.615000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.140000  1.105000  6.310000 1.275000 ;
      RECT  6.140000  1.785000  6.310000 1.955000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.900000  1.445000  9.070000 1.615000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 0.735000 0.840000 0.780000 ;
      RECT 0.550000 0.780000 3.130000 0.920000 ;
      RECT 0.550000 0.920000 0.840000 0.965000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 6.370000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.400000 1.755000 2.690000 1.800000 ;
      RECT 2.400000 1.940000 2.690000 1.985000 ;
      RECT 2.840000 0.735000 3.130000 0.780000 ;
      RECT 2.840000 0.920000 3.130000 0.965000 ;
      RECT 2.935000 0.965000 3.130000 1.120000 ;
      RECT 2.935000 1.120000 6.370000 1.260000 ;
      RECT 5.620000 1.415000 5.910000 1.460000 ;
      RECT 5.620000 1.460000 9.130000 1.600000 ;
      RECT 5.620000 1.600000 5.910000 1.645000 ;
      RECT 6.080000 1.075000 6.370000 1.120000 ;
      RECT 6.080000 1.260000 6.370000 1.305000 ;
      RECT 6.080000 1.755000 6.370000 1.800000 ;
      RECT 6.080000 1.940000 6.370000 1.985000 ;
      RECT 8.840000 1.415000 9.130000 1.460000 ;
      RECT 8.840000 1.600000 9.130000 1.645000 ;
  END
END sky130_fd_sc_hd__dfbbn_2
MACRO sky130_fd_sc_hd__dfbbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfbbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.745000 1.005000 2.155000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.615000 0.255000 11.875000 0.825000 ;
        RECT 11.615000 1.455000 11.875000 2.465000 ;
        RECT 11.665000 0.825000 11.875000 1.455000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.200000 0.255000 10.485000 0.715000 ;
        RECT 10.200000 1.630000 10.485000 2.465000 ;
        RECT 10.305000 0.715000 10.485000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.235000 1.095000 9.690000 1.325000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.585000 0.735000 3.995000 0.965000 ;
        RECT 3.585000 0.965000 3.915000 1.065000 ;
      LAYER mcon ;
        RECT 3.825000 0.765000 3.995000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.280000 0.735000 7.825000 1.065000 ;
      LAYER mcon ;
        RECT 7.575000 0.765000 7.745000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765000 0.735000 4.055000 0.780000 ;
        RECT 3.765000 0.780000 7.805000 0.920000 ;
        RECT 3.765000 0.920000 4.055000 0.965000 ;
        RECT 7.515000 0.735000 7.805000 0.780000 ;
        RECT 7.515000 0.920000 7.805000 0.965000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.840000 0.805000 ;
      RECT  0.175000  1.795000  0.840000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.235000 2.465000 ;
      RECT  1.405000  0.635000  2.125000 0.825000 ;
      RECT  1.405000  0.825000  1.575000 1.795000 ;
      RECT  1.405000  1.795000  2.125000 1.965000 ;
      RECT  1.430000  0.085000  1.785000 0.465000 ;
      RECT  1.430000  2.135000  1.785000 2.635000 ;
      RECT  1.955000  0.305000  2.125000 0.635000 ;
      RECT  1.955000  1.965000  2.125000 2.465000 ;
      RECT  2.325000  0.705000  2.545000 1.575000 ;
      RECT  2.325000  1.575000  2.825000 1.955000 ;
      RECT  2.335000  2.250000  3.165000 2.420000 ;
      RECT  2.400000  0.265000  3.415000 0.465000 ;
      RECT  2.725000  0.645000  3.075000 1.015000 ;
      RECT  2.995000  1.195000  3.415000 1.235000 ;
      RECT  2.995000  1.235000  4.345000 1.405000 ;
      RECT  2.995000  1.405000  3.165000 2.250000 ;
      RECT  3.245000  0.465000  3.415000 1.195000 ;
      RECT  3.335000  1.575000  3.585000 1.785000 ;
      RECT  3.335000  1.785000  4.685000 2.035000 ;
      RECT  3.405000  2.205000  3.785000 2.635000 ;
      RECT  3.585000  0.085000  3.755000 0.525000 ;
      RECT  3.925000  0.255000  5.075000 0.425000 ;
      RECT  3.925000  0.425000  4.255000 0.505000 ;
      RECT  4.085000  2.035000  4.255000 2.375000 ;
      RECT  4.095000  1.405000  4.345000 1.485000 ;
      RECT  4.125000  1.155000  4.345000 1.235000 ;
      RECT  4.405000  0.595000  4.735000 0.765000 ;
      RECT  4.515000  0.765000  4.735000 0.895000 ;
      RECT  4.515000  0.895000  5.825000 1.065000 ;
      RECT  4.515000  1.065000  4.685000 1.785000 ;
      RECT  4.855000  1.235000  5.185000 1.415000 ;
      RECT  4.855000  1.415000  5.860000 1.655000 ;
      RECT  4.875000  1.915000  5.205000 2.635000 ;
      RECT  4.905000  0.425000  5.075000 0.715000 ;
      RECT  5.325000  0.085000  5.675000 0.465000 ;
      RECT  5.495000  1.065000  5.825000 1.235000 ;
      RECT  6.060000  1.575000  6.295000 1.985000 ;
      RECT  6.065000  1.060000  6.405000 1.125000 ;
      RECT  6.065000  1.125000  6.740000 1.305000 ;
      RECT  6.185000  0.705000  6.405000 1.060000 ;
      RECT  6.250000  2.250000  7.080000 2.420000 ;
      RECT  6.300000  0.265000  7.080000 0.465000 ;
      RECT  6.535000  1.305000  6.740000 1.905000 ;
      RECT  6.910000  0.465000  7.080000 1.235000 ;
      RECT  6.910000  1.235000  8.260000 1.405000 ;
      RECT  6.910000  1.405000  7.080000 2.250000 ;
      RECT  7.250000  0.085000  7.575000 0.525000 ;
      RECT  7.250000  1.575000  7.500000 1.915000 ;
      RECT  7.250000  1.915000 10.030000 2.085000 ;
      RECT  7.320000  2.255000  7.700000 2.635000 ;
      RECT  7.745000  0.255000  8.955000 0.425000 ;
      RECT  7.745000  0.425000  8.075000 0.545000 ;
      RECT  7.940000  2.085000  8.110000 2.375000 ;
      RECT  8.040000  1.075000  8.260000 1.235000 ;
      RECT  8.215000  0.665000  8.615000 0.835000 ;
      RECT  8.430000  0.835000  8.615000 0.840000 ;
      RECT  8.430000  0.840000  8.600000 1.915000 ;
      RECT  8.640000  2.255000 10.030000 2.635000 ;
      RECT  8.770000  1.110000  9.055000 1.575000 ;
      RECT  8.770000  1.575000  9.555000 1.745000 ;
      RECT  8.785000  0.425000  8.955000 0.585000 ;
      RECT  8.835000  0.755000  9.475000 0.925000 ;
      RECT  8.835000  0.925000  9.055000 1.110000 ;
      RECT  9.265000  0.265000  9.475000 0.755000 ;
      RECT  9.725000  0.085000 10.030000 0.805000 ;
      RECT  9.860000  0.995000 10.125000 1.325000 ;
      RECT  9.860000  1.325000 10.030000 1.915000 ;
      RECT 10.660000  0.255000 10.975000 0.995000 ;
      RECT 10.660000  0.995000 11.495000 1.325000 ;
      RECT 10.660000  1.325000 10.975000 2.415000 ;
      RECT 11.150000  0.085000 11.445000 0.545000 ;
      RECT 11.155000  1.765000 11.445000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.610000  0.765000  0.780000 0.935000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  1.785000  1.235000 1.955000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.785000  2.615000 1.955000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  0.765000  3.075000 0.935000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  1.445000  5.835000 1.615000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  1.105000  6.295000 1.275000 ;
      RECT  6.125000  1.785000  6.295000 1.955000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.855000  1.445000  9.025000 1.615000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 0.735000 0.840000 0.780000 ;
      RECT 0.550000 0.780000 3.135000 0.920000 ;
      RECT 0.550000 0.920000 0.840000 0.965000 ;
      RECT 1.005000 1.755000 1.295000 1.800000 ;
      RECT 1.005000 1.800000 6.355000 1.940000 ;
      RECT 1.005000 1.940000 1.295000 1.985000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.845000 0.735000 3.135000 0.780000 ;
      RECT 2.845000 0.920000 3.135000 0.965000 ;
      RECT 2.920000 0.965000 3.135000 1.120000 ;
      RECT 2.920000 1.120000 6.355000 1.260000 ;
      RECT 5.605000 1.415000 5.895000 1.460000 ;
      RECT 5.605000 1.460000 9.085000 1.600000 ;
      RECT 5.605000 1.600000 5.895000 1.645000 ;
      RECT 6.065000 1.075000 6.355000 1.120000 ;
      RECT 6.065000 1.260000 6.355000 1.305000 ;
      RECT 6.065000 1.755000 6.355000 1.800000 ;
      RECT 6.065000 1.940000 6.355000 1.985000 ;
      RECT 8.795000 1.415000 9.085000 1.460000 ;
      RECT 8.795000 1.600000 9.085000 1.645000 ;
  END
END sky130_fd_sc_hd__dfbbn_1
MACRO sky130_fd_sc_hd__o21ba_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.100000 1.075000 3.595000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.075000 2.930000 1.285000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.325000 ;
        RECT 0.595000 1.325000 0.775000 1.695000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.255000 1.240000 0.595000 ;
        RECT 0.945000 0.595000 1.115000 1.495000 ;
        RECT 0.945000 1.495000 1.350000 1.695000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.430000 0.345000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 0.395000 1.865000 ;
      RECT 0.085000  1.865000 1.935000 2.035000 ;
      RECT 0.520000  2.205000 0.910000 2.635000 ;
      RECT 0.595000  0.085000 0.775000 0.825000 ;
      RECT 1.285000  0.890000 1.595000 1.060000 ;
      RECT 1.285000  1.060000 1.455000 1.325000 ;
      RECT 1.410000  0.085000 1.770000 0.485000 ;
      RECT 1.415000  2.205000 2.230000 2.635000 ;
      RECT 1.425000  0.655000 2.275000 0.825000 ;
      RECT 1.425000  0.825000 1.595000 0.890000 ;
      RECT 1.765000  0.995000 1.935000 1.865000 ;
      RECT 1.940000  0.255000 2.275000 0.655000 ;
      RECT 2.105000  0.825000 2.275000 1.455000 ;
      RECT 2.105000  1.455000 2.725000 2.035000 ;
      RECT 2.400000  2.035000 2.725000 2.465000 ;
      RECT 2.445000  0.365000 2.745000 0.735000 ;
      RECT 2.445000  0.735000 3.590000 0.905000 ;
      RECT 2.915000  0.085000 3.085000 0.555000 ;
      RECT 3.200000  1.875000 3.530000 2.635000 ;
      RECT 3.255000  0.270000 3.590000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ba_2
MACRO sky130_fd_sc_hd__o21ba_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.990000 1.075000 5.895000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.780000 1.075000 4.820000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 0.885000 1.285000 ;
        RECT 0.605000 1.285000 0.885000 1.705000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 0.255000 1.385000 0.725000 ;
        RECT 1.055000 0.725000 2.225000 0.905000 ;
        RECT 1.055000 0.905000 1.455000 1.445000 ;
        RECT 1.055000 1.445000 2.225000 1.705000 ;
        RECT 1.895000 0.255000 2.225000 0.725000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.265000 0.545000 0.855000 ;
      RECT 0.085000  0.855000 0.255000 1.455000 ;
      RECT 0.085000  1.455000 0.435000 1.875000 ;
      RECT 0.085000  1.875000 2.565000 2.045000 ;
      RECT 0.085000  2.045000 0.435000 2.465000 ;
      RECT 0.635000  2.215000 0.965000 2.635000 ;
      RECT 0.715000  0.085000 0.885000 0.905000 ;
      RECT 1.475000  2.215000 1.805000 2.635000 ;
      RECT 1.555000  0.085000 1.725000 0.555000 ;
      RECT 1.625000  1.075000 2.565000 1.275000 ;
      RECT 2.315000  2.215000 2.645000 2.635000 ;
      RECT 2.395000  0.085000 2.565000 0.555000 ;
      RECT 2.395000  0.725000 3.585000 0.895000 ;
      RECT 2.395000  0.895000 2.565000 1.075000 ;
      RECT 2.395000  1.445000 2.905000 1.615000 ;
      RECT 2.395000  1.615000 2.565000 1.875000 ;
      RECT 2.735000  1.075000 3.135000 1.245000 ;
      RECT 2.735000  1.245000 2.905000 1.445000 ;
      RECT 2.805000  0.255000 4.005000 0.475000 ;
      RECT 2.815000  1.795000 4.380000 1.965000 ;
      RECT 2.815000  1.965000 2.985000 2.465000 ;
      RECT 3.200000  2.135000 3.450000 2.635000 ;
      RECT 3.235000  0.645000 3.585000 0.725000 ;
      RECT 3.395000  0.895000 3.585000 1.795000 ;
      RECT 3.685000  2.135000 3.925000 2.295000 ;
      RECT 3.685000  2.295000 4.765000 2.465000 ;
      RECT 3.755000  0.475000 4.005000 0.725000 ;
      RECT 3.755000  0.725000 5.710000 0.905000 ;
      RECT 4.135000  1.445000 4.380000 1.795000 ;
      RECT 4.135000  1.965000 4.380000 2.125000 ;
      RECT 4.175000  0.085000 4.345000 0.555000 ;
      RECT 4.515000  0.255000 4.845000 0.725000 ;
      RECT 4.595000  1.455000 5.710000 1.665000 ;
      RECT 4.595000  1.665000 4.765000 2.295000 ;
      RECT 4.935000  1.835000 5.265000 2.635000 ;
      RECT 5.015000  0.085000 5.185000 0.555000 ;
      RECT 5.355000  0.265000 5.710000 0.725000 ;
      RECT 5.435000  1.665000 5.710000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ba_4
MACRO sky130_fd_sc_hd__o21ba_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.950000 1.075000 3.595000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.075000 2.780000 1.285000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 0.995000 1.360000 1.325000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.450000 0.445000 0.825000 ;
        RECT 0.085000 0.825000 0.340000 1.480000 ;
        RECT 0.085000 1.480000 0.425000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.510000  0.995000 0.860000 1.325000 ;
      RECT 0.595000  1.325000 0.860000 1.865000 ;
      RECT 0.595000  1.865000 2.575000 2.035000 ;
      RECT 0.595000  2.205000 1.005000 2.635000 ;
      RECT 0.710000  0.085000 0.880000 0.825000 ;
      RECT 1.075000  1.525000 1.700000 1.695000 ;
      RECT 1.160000  0.450000 1.330000 0.655000 ;
      RECT 1.160000  0.655000 1.700000 0.825000 ;
      RECT 1.530000  0.825000 1.700000 1.525000 ;
      RECT 1.750000  2.215000 2.080000 2.635000 ;
      RECT 1.870000  0.255000 2.040000 1.455000 ;
      RECT 1.870000  1.455000 2.575000 1.865000 ;
      RECT 2.250000  2.035000 2.575000 2.465000 ;
      RECT 2.270000  0.255000 2.600000 0.735000 ;
      RECT 2.270000  0.735000 3.440000 0.905000 ;
      RECT 2.770000  0.085000 2.940000 0.555000 ;
      RECT 3.050000  1.535000 3.380000 2.635000 ;
      RECT 3.110000  0.270000 3.440000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ba_1
MACRO sky130_fd_sc_hd__nor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 0.655000 1.755000 1.665000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.995000 0.975000 1.325000 ;
        RECT 0.595000 1.325000 0.830000 2.005000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.425000 1.325000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.604500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.385000 0.345000 0.655000 ;
        RECT 0.090000 0.655000 1.315000 0.825000 ;
        RECT 0.090000 1.495000 0.425000 2.280000 ;
        RECT 0.090000 2.280000 1.170000 2.450000 ;
        RECT 1.000000 1.495000 1.315000 1.665000 ;
        RECT 1.000000 1.665000 1.170000 2.280000 ;
        RECT 1.015000 0.385000 1.185000 0.655000 ;
        RECT 1.145000 0.825000 1.315000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 1.355000  0.085000 1.685000 0.485000 ;
      RECT 1.435000  1.835000 1.750000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__nor3_1
MACRO sky130_fd_sc_hd__nor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 1.075000 0.965000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135000 1.075000 2.185000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 1.075000 2.965000 1.285000 ;
        RECT 2.375000 1.285000 2.640000 1.625000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 3.595000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.755000 0.255000 3.085000 0.725000 ;
        RECT 2.835000 1.455000 3.595000 1.625000 ;
        RECT 2.835000 1.625000 3.045000 2.125000 ;
        RECT 3.135000 0.905000 3.595000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.150000  1.455000 2.085000 1.625000 ;
      RECT 0.150000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.995000  1.625000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.795000 1.665000 2.295000 ;
      RECT 1.415000  2.295000 3.465000 2.465000 ;
      RECT 1.835000  1.625000 2.085000 2.125000 ;
      RECT 1.875000  0.085000 2.585000 0.555000 ;
      RECT 2.415000  1.795000 2.625000 2.295000 ;
      RECT 3.215000  1.795000 3.465000 2.295000 ;
      RECT 3.255000  0.085000 3.545000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__nor3_2
MACRO sky130_fd_sc_hd__nor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.825000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095000 1.075000 3.685000 1.285000 ;
        RECT 3.515000 1.285000 3.685000 1.445000 ;
        RECT 3.515000 1.445000 5.165000 1.615000 ;
        RECT 4.995000 1.075000 5.415000 1.285000 ;
        RECT 4.995000 1.285000 5.165000 1.445000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.855000 1.075000 4.765000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 5.895000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 3.515000 1.785000 5.895000 1.955000 ;
        RECT 3.515000 1.955000 4.605000 1.965000 ;
        RECT 3.515000 1.965000 3.765000 2.125000 ;
        RECT 3.895000 0.255000 4.225000 0.725000 ;
        RECT 4.355000 1.965000 4.605000 2.125000 ;
        RECT 4.735000 0.255000 5.065000 0.725000 ;
        RECT 5.605000 0.255000 5.895000 0.725000 ;
        RECT 5.605000 0.905000 5.895000 1.785000 ;
        RECT 5.615000 1.955000 5.895000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.150000  1.455000 2.085000 1.625000 ;
      RECT 0.150000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.995000  1.625000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.795000 1.665000 2.635000 ;
      RECT 1.835000  1.625000 2.085000 2.085000 ;
      RECT 1.835000  2.085000 2.925000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.255000  1.455000 3.345000 1.625000 ;
      RECT 2.255000  1.625000 2.505000 1.915000 ;
      RECT 2.675000  1.795000 2.925000 2.085000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 3.095000  1.625000 3.345000 2.295000 ;
      RECT 3.095000  2.295000 5.025000 2.465000 ;
      RECT 3.555000  0.085000 3.725000 0.555000 ;
      RECT 3.935000  2.135000 4.185000 2.295000 ;
      RECT 4.395000  0.085000 4.565000 0.555000 ;
      RECT 4.775000  2.135000 5.025000 2.295000 ;
      RECT 5.195000  2.125000 5.445000 2.465000 ;
      RECT 5.235000  0.085000 5.405000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.125000 2.615000 2.295000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.125000 5.375000 2.295000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 2.385000 2.065000 2.680000 2.140000 ;
      RECT 2.385000 2.140000 5.440000 2.280000 ;
      RECT 2.385000 2.280000 2.680000 2.335000 ;
      RECT 5.145000 2.065000 5.440000 2.140000 ;
      RECT 5.145000 2.280000 5.440000 2.335000 ;
  END
END sky130_fd_sc_hd__nor3_4
MACRO sky130_fd_sc_hd__or3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.995000 1.430000 1.325000 ;
        RECT 0.605000 1.325000 0.830000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 2.125000 1.280000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.435000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 0.415000 2.215000 0.760000 ;
        RECT 1.940000 1.495000 2.215000 2.465000 ;
        RECT 2.045000 0.760000 2.215000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.105000  0.305000 0.360000 0.655000 ;
      RECT 0.105000  0.655000 1.770000 0.825000 ;
      RECT 0.105000  1.495000 0.435000 1.785000 ;
      RECT 0.105000  1.785000 1.270000 1.955000 ;
      RECT 0.530000  0.085000 0.860000 0.485000 ;
      RECT 1.030000  0.305000 1.200000 0.655000 ;
      RECT 1.100000  1.495000 1.770000 1.665000 ;
      RECT 1.100000  1.665000 1.270000 1.785000 ;
      RECT 1.370000  0.085000 1.750000 0.485000 ;
      RECT 1.450000  1.835000 1.730000 2.635000 ;
      RECT 1.600000  0.825000 1.770000 0.995000 ;
      RECT 1.600000  0.995000 1.875000 1.325000 ;
      RECT 1.600000  1.325000 1.770000 1.495000 ;
      RECT 2.385000  0.085000 2.675000 0.915000 ;
      RECT 2.385000  1.430000 2.675000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__or3_2
MACRO sky130_fd_sc_hd__or3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.600000 0.995000 1.425000 1.325000 ;
        RECT 0.600000 1.325000 0.795000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 2.125000 1.275000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.430000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.415000 2.210000 0.760000 ;
        RECT 1.935000 1.495000 2.210000 2.465000 ;
        RECT 2.040000 0.760000 2.210000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.100000  0.305000 0.355000 0.655000 ;
      RECT 0.100000  0.655000 1.765000 0.825000 ;
      RECT 0.105000  1.495000 0.430000 1.785000 ;
      RECT 0.105000  1.785000 1.275000 1.955000 ;
      RECT 0.525000  0.085000 0.855000 0.485000 ;
      RECT 1.025000  0.305000 1.195000 0.655000 ;
      RECT 1.105000  1.495000 1.765000 1.665000 ;
      RECT 1.105000  1.665000 1.275000 1.785000 ;
      RECT 1.365000  0.085000 1.745000 0.485000 ;
      RECT 1.445000  1.835000 1.725000 2.635000 ;
      RECT 1.595000  0.825000 1.765000 0.995000 ;
      RECT 1.595000  0.995000 1.870000 1.325000 ;
      RECT 1.595000  1.325000 1.765000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__or3_1
MACRO sky130_fd_sc_hd__or3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 1.075000 1.700000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 1.075000 1.055000 1.325000 ;
        RECT 0.595000 1.325000 0.830000 2.050000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.305000 0.265000 2.635000 0.735000 ;
        RECT 2.305000 0.735000 4.055000 0.905000 ;
        RECT 2.345000 1.455000 4.055000 1.625000 ;
        RECT 2.345000 1.625000 2.595000 2.465000 ;
        RECT 3.145000 0.265000 3.475000 0.735000 ;
        RECT 3.185000 1.625000 3.435000 2.465000 ;
        RECT 3.765000 0.905000 4.055000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.255000 0.425000 0.725000 ;
      RECT 0.085000  0.725000 2.090000 0.905000 ;
      RECT 0.085000  1.495000 0.425000 2.295000 ;
      RECT 0.085000  2.295000 1.265000 2.465000 ;
      RECT 0.595000  0.085000 0.765000 0.555000 ;
      RECT 0.935000  0.255000 1.265000 0.725000 ;
      RECT 1.000000  1.495000 2.090000 1.665000 ;
      RECT 1.000000  1.665000 1.265000 2.295000 ;
      RECT 1.435000  0.085000 2.135000 0.555000 ;
      RECT 1.435000  1.835000 2.135000 2.635000 ;
      RECT 1.870000  0.905000 2.090000 1.075000 ;
      RECT 1.870000  1.075000 3.595000 1.245000 ;
      RECT 1.870000  1.245000 2.090000 1.495000 ;
      RECT 2.765000  1.795000 3.015000 2.635000 ;
      RECT 2.805000  0.085000 2.975000 0.555000 ;
      RECT 3.605000  1.795000 3.855000 2.635000 ;
      RECT 3.645000  0.085000 3.815000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__or3_4
MACRO sky130_fd_sc_hd__lpflow_inputiso0n_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso0n_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 0.775000 1.325000 ;
        RECT 0.100000 1.325000 0.365000 1.685000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.075000 1.335000 1.325000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.657000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655000 0.255000 2.215000 0.545000 ;
        RECT 1.755000 1.915000 2.215000 2.465000 ;
        RECT 1.965000 0.545000 2.215000 1.915000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.285000  0.355000 0.615000 0.715000 ;
      RECT 0.285000  0.715000 1.675000 0.905000 ;
      RECT 0.285000  1.965000 0.565000 2.635000 ;
      RECT 0.735000  1.575000 1.675000 1.745000 ;
      RECT 0.735000  1.745000 1.035000 2.295000 ;
      RECT 1.235000  0.085000 1.485000 0.545000 ;
      RECT 1.235000  1.915000 1.565000 2.635000 ;
      RECT 1.505000  0.905000 1.675000 0.995000 ;
      RECT 1.505000  0.995000 1.795000 1.325000 ;
      RECT 1.505000  1.325000 1.675000 1.575000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso0n_1
MACRO sky130_fd_sc_hd__tapvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvgnd_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.315000 0.845000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.085000 2.095000 0.375000 2.325000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  1.470000 0.375000 2.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.125000 0.315000 2.295000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__tapvgnd_1
MACRO sky130_fd_sc_hd__and4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.625000 0.775000 1.955000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.765000 0.815000 0.945000 ;
        RECT 0.605000 0.945000 1.225000 1.115000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895000 0.415000 3.080000 0.995000 ;
        RECT 2.895000 0.995000 3.125000 1.325000 ;
        RECT 2.895000 1.325000 3.080000 1.635000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 0.420000 3.545000 0.995000 ;
        RECT 3.350000 0.995000 3.605000 1.325000 ;
        RECT 3.350000 1.325000 3.545000 1.635000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.425400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.255000 0.255000 4.515000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.285000 ;
      RECT 0.085000  1.285000 1.215000 1.455000 ;
      RECT 0.085000  1.455000 0.255000 2.135000 ;
      RECT 0.085000  2.135000 0.345000 2.465000 ;
      RECT 0.655000  0.085000 0.985000 0.465000 ;
      RECT 0.655000  2.255000 0.985000 2.635000 ;
      RECT 1.045000  1.455000 1.215000 1.575000 ;
      RECT 1.045000  1.575000 1.625000 1.745000 ;
      RECT 1.165000  0.255000 2.645000 0.425000 ;
      RECT 1.165000  0.425000 1.565000 0.755000 ;
      RECT 1.225000  1.915000 1.965000 2.085000 ;
      RECT 1.225000  2.085000 1.415000 2.465000 ;
      RECT 1.395000  0.755000 1.565000 1.235000 ;
      RECT 1.395000  1.235000 1.965000 1.405000 ;
      RECT 1.665000  2.255000 1.995000 2.635000 ;
      RECT 1.755000  0.595000 2.305000 0.925000 ;
      RECT 1.795000  1.405000 1.965000 1.915000 ;
      RECT 2.135000  0.925000 2.305000 1.915000 ;
      RECT 2.135000  1.915000 4.085000 2.085000 ;
      RECT 2.205000  2.085000 2.375000 2.465000 ;
      RECT 2.475000  0.425000 2.645000 1.325000 ;
      RECT 2.570000  2.255000 2.900000 2.635000 ;
      RECT 3.160000  2.085000 3.330000 2.465000 ;
      RECT 3.755000  0.085000 4.085000 0.465000 ;
      RECT 3.755000  2.255000 4.085000 2.635000 ;
      RECT 3.915000  0.995000 4.085000 1.915000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__and4bb_1
MACRO sky130_fd_sc_hd__and4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.485000 0.995000 5.845000 1.620000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.765000 0.780000 1.635000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.250000 0.755000 3.545000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.680000 0.995000 3.080000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 0.650000 2.080000 0.820000 ;
        RECT 0.960000 0.820000 1.240000 1.545000 ;
        RECT 0.960000 1.545000 2.160000 1.715000 ;
        RECT 1.070000 0.255000 1.240000 0.650000 ;
        RECT 1.910000 0.255000 2.080000 0.650000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.260000 1.915000 ;
      RECT 0.085000  1.915000 4.490000 2.085000 ;
      RECT 0.085000  2.085000 0.345000 2.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 0.570000  0.085000 0.900000 0.470000 ;
      RECT 1.410000  0.085000 1.740000 0.470000 ;
      RECT 1.410000  1.075000 2.500000 1.245000 ;
      RECT 1.410000  2.255000 1.740000 2.635000 ;
      RECT 2.250000  2.255000 2.580000 2.635000 ;
      RECT 2.270000  0.085000 2.600000 0.445000 ;
      RECT 2.330000  0.615000 2.940000 0.785000 ;
      RECT 2.330000  0.785000 2.500000 1.075000 ;
      RECT 2.330000  1.245000 2.500000 1.545000 ;
      RECT 2.330000  1.545000 4.150000 1.715000 ;
      RECT 2.770000  0.300000 4.610000 0.470000 ;
      RECT 2.770000  0.470000 2.940000 0.615000 ;
      RECT 3.330000  2.255000 3.660000 2.635000 ;
      RECT 3.730000  0.995000 3.900000 1.155000 ;
      RECT 3.730000  1.155000 4.490000 1.325000 ;
      RECT 4.255000  0.470000 4.610000 0.810000 ;
      RECT 4.320000  1.325000 4.490000 1.915000 ;
      RECT 4.360000  2.255000 5.370000 2.635000 ;
      RECT 4.950000  0.655000 5.805000 0.825000 ;
      RECT 4.950000  0.825000 5.120000 1.915000 ;
      RECT 4.950000  1.915000 5.805000 2.085000 ;
      RECT 4.975000  0.085000 5.305000 0.465000 ;
      RECT 5.635000  0.255000 5.805000 0.655000 ;
      RECT 5.635000  2.085000 5.805000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__and4bb_4
MACRO sky130_fd_sc_hd__and4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.995000 0.330000 1.635000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 0.765000 4.175000 1.305000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.910000 0.420000 3.175000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 0.425000 3.655000 1.405000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.990000 1.545000 1.320000 1.715000 ;
        RECT 1.015000 0.255000 1.240000 1.545000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.670000 0.805000 ;
      RECT 0.175000  1.885000 1.925000 2.055000 ;
      RECT 0.175000  2.055000 0.345000 2.465000 ;
      RECT 0.500000  0.805000 0.670000 1.885000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 1.410000  0.085000 1.740000 0.465000 ;
      RECT 1.415000  0.635000 2.405000 0.805000 ;
      RECT 1.415000  0.805000 1.585000 1.325000 ;
      RECT 1.490000  2.255000 2.160000 2.635000 ;
      RECT 1.755000  0.995000 2.065000 1.325000 ;
      RECT 1.755000  1.325000 1.925000 1.885000 ;
      RECT 2.010000  0.255000 2.180000 0.635000 ;
      RECT 2.235000  0.805000 2.405000 1.915000 ;
      RECT 2.235000  1.915000 3.415000 2.085000 ;
      RECT 2.395000  2.085000 2.565000 2.465000 ;
      RECT 2.575000  1.400000 2.745000 1.575000 ;
      RECT 2.575000  1.575000 3.755000 1.745000 ;
      RECT 2.735000  2.255000 3.075000 2.635000 ;
      RECT 3.245000  2.085000 3.415000 2.465000 ;
      RECT 3.585000  1.745000 3.755000 1.915000 ;
      RECT 3.585000  1.915000 4.515000 2.085000 ;
      RECT 3.755000  2.255000 4.085000 2.635000 ;
      RECT 3.835000  0.085000 4.085000 0.585000 ;
      RECT 4.255000  0.255000 4.515000 0.585000 ;
      RECT 4.255000  2.085000 4.515000 2.465000 ;
      RECT 4.345000  0.585000 4.515000 1.915000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__and4bb_2
MACRO sky130_fd_sc_hd__a2bb2o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 0.995000 1.675000 1.615000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845000 0.995000 2.135000 1.375000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.730000 0.765000 3.990000 1.655000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.050000 1.355000 3.530000 1.655000 ;
        RECT 3.270000 0.765000 3.530000 1.355000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 0.255000 0.780000 0.810000 ;
        RECT 0.525000 0.810000 0.695000 1.525000 ;
        RECT 0.525000 1.525000 0.780000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125000 -0.085000 0.295000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.185000  0.085000 0.355000 0.930000 ;
      RECT 0.185000  1.445000 0.355000 2.635000 ;
      RECT 0.865000  0.995000 1.120000 1.325000 ;
      RECT 0.950000  0.085000 1.380000 0.530000 ;
      RECT 0.950000  1.325000 1.120000 1.805000 ;
      RECT 0.950000  1.805000 1.710000 1.975000 ;
      RECT 0.950000  2.235000 1.280000 2.635000 ;
      RECT 1.540000  1.975000 1.710000 2.200000 ;
      RECT 1.540000  2.200000 2.670000 2.370000 ;
      RECT 1.615000  0.255000 1.785000 0.655000 ;
      RECT 1.615000  0.655000 2.510000 0.825000 ;
      RECT 1.955000  0.085000 2.690000 0.485000 ;
      RECT 1.975000  1.545000 2.510000 1.715000 ;
      RECT 1.975000  1.715000 2.145000 1.905000 ;
      RECT 2.340000  0.825000 2.510000 1.545000 ;
      RECT 2.440000  1.895000 2.850000 2.065000 ;
      RECT 2.440000  2.065000 2.670000 2.200000 ;
      RECT 2.500000  2.370000 2.670000 2.465000 ;
      RECT 2.680000  0.700000 3.030000 0.870000 ;
      RECT 2.680000  0.870000 2.850000 1.895000 ;
      RECT 2.860000  0.255000 3.030000 0.700000 ;
      RECT 2.875000  2.255000 3.205000 2.425000 ;
      RECT 3.035000  1.835000 3.965000 2.005000 ;
      RECT 3.035000  2.005000 3.205000 2.255000 ;
      RECT 3.375000  2.175000 3.625000 2.635000 ;
      RECT 3.605000  0.085000 4.005000 0.595000 ;
      RECT 3.795000  2.005000 3.965000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a2bb2o_2
MACRO sky130_fd_sc_hd__a2bb2o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 0.995000 1.240000 1.615000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.410000 0.995000 1.700000 1.375000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.280000 0.765000 3.540000 1.655000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.600000 1.355000 3.080000 1.655000 ;
        RECT 2.820000 0.765000 3.080000 1.355000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.345000 0.810000 ;
        RECT 0.085000 0.810000 0.260000 1.525000 ;
        RECT 0.085000 1.525000 0.345000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.430000  0.995000 0.685000 1.325000 ;
      RECT 0.515000  0.085000 0.945000 0.530000 ;
      RECT 0.515000  1.325000 0.685000 1.805000 ;
      RECT 0.515000  1.805000 1.275000 1.975000 ;
      RECT 0.515000  2.235000 0.845000 2.635000 ;
      RECT 1.105000  1.975000 1.275000 2.200000 ;
      RECT 1.105000  2.200000 2.245000 2.370000 ;
      RECT 1.180000  0.255000 1.350000 0.655000 ;
      RECT 1.180000  0.655000 2.060000 0.825000 ;
      RECT 1.520000  0.085000 2.240000 0.485000 ;
      RECT 1.540000  1.545000 2.060000 1.715000 ;
      RECT 1.540000  1.715000 1.710000 1.905000 ;
      RECT 1.890000  0.825000 2.060000 1.545000 ;
      RECT 1.990000  1.895000 2.400000 2.065000 ;
      RECT 1.990000  2.065000 2.245000 2.200000 ;
      RECT 1.990000  2.370000 2.245000 2.465000 ;
      RECT 2.230000  0.700000 2.580000 0.870000 ;
      RECT 2.230000  0.870000 2.400000 1.895000 ;
      RECT 2.410000  0.255000 2.580000 0.700000 ;
      RECT 2.415000  2.255000 2.745000 2.425000 ;
      RECT 2.575000  1.835000 3.515000 2.005000 ;
      RECT 2.575000  2.005000 2.745000 2.255000 ;
      RECT 2.915000  2.175000 3.165000 2.635000 ;
      RECT 3.155000  0.085000 3.555000 0.595000 ;
      RECT 3.335000  2.005000 3.515000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a2bb2o_1
MACRO sky130_fd_sc_hd__a2bb2o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.075000 3.645000 1.325000 ;
        RECT 3.475000 1.325000 3.645000 1.445000 ;
        RECT 3.475000 1.445000 4.965000 1.615000 ;
        RECT 4.605000 1.075000 4.965000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 1.075000 4.435000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.575000 1.445000 ;
        RECT 0.085000 1.445000 1.685000 1.615000 ;
        RECT 1.515000 1.075000 1.895000 1.245000 ;
        RECT 1.515000 1.245000 1.685000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.075000 1.345000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235000 0.275000 5.565000 0.725000 ;
        RECT 5.235000 0.725000 6.920000 0.905000 ;
        RECT 5.275000 1.785000 6.365000 1.955000 ;
        RECT 5.275000 1.955000 5.525000 2.465000 ;
        RECT 6.075000 0.275000 6.405000 0.725000 ;
        RECT 6.115000 1.415000 6.920000 1.655000 ;
        RECT 6.115000 1.655000 6.365000 1.785000 ;
        RECT 6.115000 1.955000 6.365000 2.465000 ;
        RECT 6.610000 0.905000 6.920000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.135000  1.785000 2.065000 1.955000 ;
      RECT 0.135000  1.955000 0.385000 2.465000 ;
      RECT 0.175000  0.085000 0.345000 0.895000 ;
      RECT 0.515000  0.255000 1.685000 0.475000 ;
      RECT 0.515000  0.475000 0.765000 0.905000 ;
      RECT 0.555000  2.125000 0.805000 2.635000 ;
      RECT 0.935000  0.645000 1.270000 0.735000 ;
      RECT 0.935000  0.735000 2.525000 0.905000 ;
      RECT 0.975000  1.955000 1.225000 2.465000 ;
      RECT 1.395000  2.125000 1.645000 2.635000 ;
      RECT 1.815000  1.955000 2.065000 2.295000 ;
      RECT 1.815000  2.295000 2.905000 2.465000 ;
      RECT 1.855000  0.085000 2.025000 0.555000 ;
      RECT 1.855000  1.455000 2.065000 1.785000 ;
      RECT 2.195000  0.255000 2.525000 0.735000 ;
      RECT 2.235000  0.905000 2.445000 1.415000 ;
      RECT 2.235000  1.415000 2.620000 1.965000 ;
      RECT 2.235000  1.965000 2.485000 2.125000 ;
      RECT 2.615000  1.075000 3.145000 1.245000 ;
      RECT 2.655000  2.135000 2.905000 2.295000 ;
      RECT 2.695000  0.085000 3.385000 0.555000 ;
      RECT 2.955000  0.725000 4.725000 0.905000 ;
      RECT 2.955000  0.905000 3.145000 1.075000 ;
      RECT 2.955000  1.245000 3.145000 1.495000 ;
      RECT 2.955000  1.495000 3.305000 1.665000 ;
      RECT 3.135000  1.665000 3.305000 1.785000 ;
      RECT 3.135000  1.785000 4.265000 1.965000 ;
      RECT 3.175000  2.135000 3.425000 2.635000 ;
      RECT 3.555000  0.255000 3.885000 0.725000 ;
      RECT 3.595000  2.135000 3.845000 2.295000 ;
      RECT 3.595000  2.295000 4.685000 2.465000 ;
      RECT 4.015000  1.965000 4.265000 2.125000 ;
      RECT 4.055000  0.085000 4.225000 0.555000 ;
      RECT 4.395000  0.255000 4.725000 0.725000 ;
      RECT 4.435000  1.785000 4.685000 2.295000 ;
      RECT 4.855000  1.795000 5.105000 2.635000 ;
      RECT 4.895000  0.085000 5.065000 0.895000 ;
      RECT 5.135000  1.075000 6.440000 1.245000 ;
      RECT 5.135000  1.245000 5.460000 1.615000 ;
      RECT 5.695000  2.165000 5.945000 2.635000 ;
      RECT 5.735000  0.085000 5.905000 0.555000 ;
      RECT 6.535000  1.825000 6.785000 2.635000 ;
      RECT 6.575000  0.085000 6.745000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.450000  1.445000 2.620000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.230000  1.445000 5.400000 1.615000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 2.390000 1.415000 2.680000 1.460000 ;
      RECT 2.390000 1.460000 5.460000 1.600000 ;
      RECT 2.390000 1.600000 2.680000 1.645000 ;
      RECT 5.170000 1.415000 5.460000 1.460000 ;
      RECT 5.170000 1.600000 5.460000 1.645000 ;
  END
END sky130_fd_sc_hd__a2bb2o_4
MACRO sky130_fd_sc_hd__o21a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 0.995000 3.125000 1.450000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 1.025000 2.610000 1.400000 ;
        RECT 2.405000 1.400000 2.610000 1.985000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 1.010000 1.855000 1.615000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 0.255000 0.775000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  1.635000 0.345000 2.635000 ;
      RECT 0.105000  0.085000 0.345000 0.885000 ;
      RECT 0.945000  0.085000 1.275000 0.465000 ;
      RECT 0.945000  0.635000 1.795000 0.840000 ;
      RECT 0.945000  0.840000 1.275000 1.330000 ;
      RECT 0.945000  2.185000 1.795000 2.635000 ;
      RECT 1.105000  1.330000 1.275000 1.785000 ;
      RECT 1.105000  1.785000 2.225000 2.005000 ;
      RECT 1.465000  0.255000 1.795000 0.635000 ;
      RECT 1.965000  0.465000 2.175000 0.635000 ;
      RECT 1.965000  0.635000 3.120000 0.825000 ;
      RECT 1.965000  2.005000 2.225000 2.465000 ;
      RECT 2.345000  0.085000 2.675000 0.465000 ;
      RECT 2.795000  1.650000 3.120000 2.635000 ;
      RECT 2.845000  0.495000 3.120000 0.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o21a_2
MACRO sky130_fd_sc_hd__o21a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.345000 1.075000 2.675000 1.275000 ;
        RECT 2.445000 1.275000 2.675000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.705000 1.075000 2.035000 1.095000 ;
        RECT 1.705000 1.095000 2.155000 1.275000 ;
        RECT 1.940000 1.275000 2.155000 2.390000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.535000 1.305000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 1.030000 ;
        RECT 0.085000 1.030000 0.365000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.535000  1.860000 1.245000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 0.595000  0.715000 1.305000 0.905000 ;
      RECT 0.595000  0.905000 0.880000 1.475000 ;
      RECT 0.595000  1.475000 1.745000 1.690000 ;
      RECT 1.005000  0.255000 1.365000 0.520000 ;
      RECT 1.005000  0.520000 1.360000 0.525000 ;
      RECT 1.005000  0.525000 1.355000 0.535000 ;
      RECT 1.005000  0.535000 1.350000 0.540000 ;
      RECT 1.005000  0.540000 1.345000 0.550000 ;
      RECT 1.005000  0.550000 1.340000 0.555000 ;
      RECT 1.005000  0.555000 1.330000 0.565000 ;
      RECT 1.005000  0.565000 1.320000 0.575000 ;
      RECT 1.005000  0.575000 1.305000 0.715000 ;
      RECT 1.415000  1.690000 1.745000 2.465000 ;
      RECT 1.495000  0.635000 1.825000 0.715000 ;
      RECT 1.495000  0.715000 2.675000 0.905000 ;
      RECT 1.995000  0.085000 2.165000 0.545000 ;
      RECT 2.335000  0.255000 2.675000 0.715000 ;
      RECT 2.335000  1.915000 2.665000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__o21a_1
MACRO sky130_fd_sc_hd__o21a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.480000 0.990000 3.785000 1.495000 ;
        RECT 3.480000 1.495000 5.400000 1.705000 ;
        RECT 5.030000 0.995000 5.400000 1.495000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.140000 0.995000 4.690000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485000 1.075000 3.155000 1.615000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.635000 1.715000 0.805000 ;
        RECT 0.090000 0.805000 0.320000 1.530000 ;
        RECT 0.090000 1.530000 1.955000 1.700000 ;
        RECT 0.595000 0.615000 1.715000 0.635000 ;
        RECT 0.915000 1.700000 1.105000 2.465000 ;
        RECT 1.775000 1.700000 1.955000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.415000  1.870000 0.745000 2.635000 ;
      RECT 0.490000  0.995000 2.315000 1.335000 ;
      RECT 0.955000  0.085000 1.285000 0.445000 ;
      RECT 1.275000  1.870000 1.605000 2.635000 ;
      RECT 1.815000  0.085000 2.145000 0.465000 ;
      RECT 2.115000  0.655000 3.095000 0.870000 ;
      RECT 2.115000  0.870000 2.315000 0.995000 ;
      RECT 2.125000  1.335000 2.315000 1.830000 ;
      RECT 2.125000  1.830000 2.845000 1.875000 ;
      RECT 2.125000  1.875000 4.545000 2.085000 ;
      RECT 2.135000  2.255000 2.485000 2.635000 ;
      RECT 2.335000  0.255000 3.605000 0.485000 ;
      RECT 2.655000  2.085000 4.545000 2.105000 ;
      RECT 2.655000  2.105000 2.845000 2.465000 ;
      RECT 3.015000  2.275000 3.685000 2.635000 ;
      RECT 3.275000  0.485000 3.605000 0.615000 ;
      RECT 3.275000  0.615000 5.405000 0.785000 ;
      RECT 3.775000  0.085000 4.115000 0.445000 ;
      RECT 4.215000  2.105000 4.545000 2.445000 ;
      RECT 4.645000  0.085000 4.975000 0.445000 ;
      RECT 5.075000  1.935000 5.435000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__o21a_4
MACRO sky130_fd_sc_hd__dfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfstp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.005000 2.180000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.810000 1.495000 9.575000 1.615000 ;
        RECT 8.810000 1.615000 9.140000 2.460000 ;
        RECT 8.890000 0.265000 9.135000 0.765000 ;
        RECT 8.890000 0.765000 9.575000 0.825000 ;
        RECT 8.975000 0.825000 9.575000 0.855000 ;
        RECT 8.975000 1.445000 9.575000 1.495000 ;
        RECT 8.990000 0.855000 9.575000 0.895000 ;
        RECT 9.020000 0.895000 9.575000 1.445000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 0.735000 4.020000 1.065000 ;
      LAYER mcon ;
        RECT 3.825000 0.765000 3.995000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.660000 0.735000 7.340000 1.005000 ;
        RECT 6.660000 1.005000 7.010000 1.065000 ;
      LAYER mcon ;
        RECT 7.045000 0.765000 7.215000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765000 0.735000 4.055000 0.780000 ;
        RECT 3.765000 0.780000 7.275000 0.920000 ;
        RECT 3.765000 0.920000 4.055000 0.965000 ;
        RECT 6.985000 0.735000 7.275000 0.780000 ;
        RECT 6.985000 0.920000 7.275000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.835000 0.805000 ;
      RECT 0.085000  1.795000 0.835000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.605000  0.805000 0.835000 1.795000 ;
      RECT 1.005000  0.565000 1.235000 2.045000 ;
      RECT 1.015000  0.345000 1.235000 0.565000 ;
      RECT 1.015000  2.045000 1.235000 2.465000 ;
      RECT 1.430000  0.635000 2.125000 0.825000 ;
      RECT 1.430000  0.825000 1.600000 1.795000 ;
      RECT 1.430000  1.795000 2.125000 1.965000 ;
      RECT 1.455000  0.085000 1.785000 0.465000 ;
      RECT 1.455000  2.135000 1.785000 2.635000 ;
      RECT 1.955000  0.305000 2.125000 0.635000 ;
      RECT 1.955000  1.965000 2.125000 2.465000 ;
      RECT 2.350000  0.705000 2.570000 1.575000 ;
      RECT 2.350000  1.575000 2.850000 1.955000 ;
      RECT 2.360000  2.250000 3.190000 2.420000 ;
      RECT 2.425000  0.265000 3.440000 0.465000 ;
      RECT 2.750000  0.645000 3.100000 1.015000 ;
      RECT 3.020000  1.195000 3.440000 1.235000 ;
      RECT 3.020000  1.235000 4.370000 1.405000 ;
      RECT 3.020000  1.405000 3.190000 2.250000 ;
      RECT 3.270000  0.465000 3.440000 1.195000 ;
      RECT 3.360000  1.575000 3.610000 1.835000 ;
      RECT 3.360000  1.835000 4.710000 2.085000 ;
      RECT 3.430000  2.255000 3.810000 2.635000 ;
      RECT 3.610000  0.085000 4.020000 0.525000 ;
      RECT 3.990000  2.085000 4.160000 2.375000 ;
      RECT 4.120000  1.405000 4.370000 1.565000 ;
      RECT 4.310000  0.295000 4.560000 0.725000 ;
      RECT 4.310000  0.725000 4.710000 1.065000 ;
      RECT 4.330000  2.255000 4.660000 2.635000 ;
      RECT 4.540000  1.065000 4.710000 1.835000 ;
      RECT 4.760000  0.085000 5.080000 0.545000 ;
      RECT 4.880000  0.725000 6.150000 0.895000 ;
      RECT 4.880000  0.895000 5.050000 1.655000 ;
      RECT 4.880000  1.655000 5.400000 1.965000 ;
      RECT 5.110000  2.165000 5.740000 2.415000 ;
      RECT 5.220000  1.065000 5.400000 1.475000 ;
      RECT 5.570000  1.235000 7.490000 1.405000 ;
      RECT 5.570000  1.405000 5.740000 1.915000 ;
      RECT 5.570000  1.915000 6.780000 2.085000 ;
      RECT 5.570000  2.085000 5.740000 2.165000 ;
      RECT 5.640000  0.305000 6.490000 0.475000 ;
      RECT 5.800000  0.895000 6.150000 1.015000 ;
      RECT 5.910000  1.575000 7.880000 1.745000 ;
      RECT 5.920000  2.255000 6.340000 2.635000 ;
      RECT 6.320000  0.475000 6.490000 1.235000 ;
      RECT 6.540000  2.085000 6.780000 2.375000 ;
      RECT 6.690000  0.085000 7.330000 0.565000 ;
      RECT 7.010000  1.945000 7.340000 2.635000 ;
      RECT 7.140000  1.175000 7.490000 1.235000 ;
      RECT 7.510000  1.745000 7.880000 1.765000 ;
      RECT 7.510000  1.765000 7.680000 2.375000 ;
      RECT 7.530000  0.350000 7.880000 0.680000 ;
      RECT 7.690000  0.680000 7.880000 1.575000 ;
      RECT 7.970000  1.915000 8.300000 2.425000 ;
      RECT 8.050000  0.345000 8.220000 0.995000 ;
      RECT 8.050000  0.995000 8.850000 1.325000 ;
      RECT 8.050000  1.325000 8.300000 1.915000 ;
      RECT 8.390000  0.085000 8.720000 0.825000 ;
      RECT 8.470000  1.495000 8.640000 2.635000 ;
      RECT 9.305000  0.085000 9.575000 0.595000 ;
      RECT 9.310000  1.785000 9.575000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  1.785000 0.775000 1.955000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  0.765000 1.235000 0.935000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.785000 2.615000 1.955000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  0.765000 3.075000 0.935000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  1.785000 5.375000 1.955000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.225000  1.105000 5.395000 1.275000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.545000 1.755000 0.835000 1.800000 ;
      RECT 0.545000 1.800000 5.435000 1.940000 ;
      RECT 0.545000 1.940000 0.835000 1.985000 ;
      RECT 1.005000 0.735000 1.295000 0.780000 ;
      RECT 1.005000 0.780000 3.135000 0.920000 ;
      RECT 1.005000 0.920000 1.295000 0.965000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.845000 0.735000 3.135000 0.780000 ;
      RECT 2.845000 0.920000 3.135000 0.965000 ;
      RECT 2.920000 0.965000 3.135000 1.120000 ;
      RECT 2.920000 1.120000 5.455000 1.260000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 5.165000 1.075000 5.455000 1.120000 ;
      RECT 5.165000 1.260000 5.455000 1.305000 ;
  END
END sky130_fd_sc_hd__dfstp_2
MACRO sky130_fd_sc_hd__dfstp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfstp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.005000 2.180000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.320000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  8.925000 0.265000  9.170000 0.715000 ;
        RECT  8.925000 0.715000 10.955000 0.885000 ;
        RECT  8.925000 1.470000 10.955000 1.640000 ;
        RECT  8.925000 1.640000  9.170000 2.465000 ;
        RECT  9.765000 0.265000  9.935000 0.715000 ;
        RECT  9.765000 1.640000  9.935000 2.465000 ;
        RECT 10.605000 0.265000 10.955000 0.715000 ;
        RECT 10.605000 1.640000 10.955000 2.465000 ;
        RECT 10.725000 0.885000 10.955000 1.470000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 0.735000 4.020000 1.065000 ;
      LAYER mcon ;
        RECT 3.825000 0.765000 3.995000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.660000 0.735000 7.320000 1.005000 ;
        RECT 6.660000 1.005000 6.990000 1.065000 ;
      LAYER mcon ;
        RECT 7.045000 0.765000 7.215000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765000 0.735000 4.055000 0.780000 ;
        RECT 3.765000 0.780000 7.275000 0.920000 ;
        RECT 3.765000 0.920000 4.055000 0.965000 ;
        RECT 6.985000 0.735000 7.275000 0.780000 ;
        RECT 6.985000 0.920000 7.275000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.840000 0.805000 ;
      RECT  0.175000  1.795000  0.840000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.240000 2.465000 ;
      RECT  1.430000  0.635000  2.125000 0.825000 ;
      RECT  1.430000  0.825000  1.600000 1.795000 ;
      RECT  1.430000  1.795000  2.125000 1.965000 ;
      RECT  1.455000  0.085000  1.785000 0.465000 ;
      RECT  1.455000  2.135000  1.785000 2.635000 ;
      RECT  1.955000  0.305000  2.125000 0.635000 ;
      RECT  1.955000  1.965000  2.125000 2.465000 ;
      RECT  2.350000  0.705000  2.570000 1.575000 ;
      RECT  2.350000  1.575000  2.850000 1.955000 ;
      RECT  2.360000  2.250000  3.190000 2.420000 ;
      RECT  2.425000  0.265000  3.440000 0.465000 ;
      RECT  2.750000  0.645000  3.100000 1.015000 ;
      RECT  3.020000  1.195000  3.440000 1.235000 ;
      RECT  3.020000  1.235000  4.370000 1.405000 ;
      RECT  3.020000  1.405000  3.190000 2.250000 ;
      RECT  3.270000  0.465000  3.440000 1.195000 ;
      RECT  3.360000  1.575000  3.610000 1.835000 ;
      RECT  3.360000  1.835000  4.710000 2.085000 ;
      RECT  3.430000  2.255000  3.810000 2.635000 ;
      RECT  3.610000  0.085000  4.020000 0.525000 ;
      RECT  3.990000  2.085000  4.160000 2.375000 ;
      RECT  4.120000  1.405000  4.370000 1.565000 ;
      RECT  4.310000  0.295000  4.560000 0.725000 ;
      RECT  4.310000  0.725000  4.710000 1.065000 ;
      RECT  4.330000  2.255000  4.660000 2.635000 ;
      RECT  4.540000  1.065000  4.710000 1.835000 ;
      RECT  4.740000  0.085000  5.080000 0.545000 ;
      RECT  4.880000  0.725000  6.150000 0.895000 ;
      RECT  4.880000  0.895000  5.050000 1.655000 ;
      RECT  4.880000  1.655000  5.400000 1.965000 ;
      RECT  5.110000  2.165000  5.740000 2.415000 ;
      RECT  5.220000  1.065000  5.400000 1.475000 ;
      RECT  5.570000  1.235000  7.470000 1.405000 ;
      RECT  5.570000  1.405000  5.740000 1.915000 ;
      RECT  5.570000  1.915000  6.780000 2.085000 ;
      RECT  5.570000  2.085000  5.740000 2.165000 ;
      RECT  5.640000  0.305000  6.490000 0.475000 ;
      RECT  5.820000  0.895000  6.150000 1.015000 ;
      RECT  5.910000  1.575000  7.850000 1.745000 ;
      RECT  5.920000  2.255000  6.340000 2.635000 ;
      RECT  6.320000  0.475000  6.490000 1.235000 ;
      RECT  6.540000  2.085000  6.780000 2.375000 ;
      RECT  6.670000  0.085000  7.330000 0.565000 ;
      RECT  7.010000  1.945000  7.340000 2.635000 ;
      RECT  7.140000  1.175000  7.470000 1.235000 ;
      RECT  7.510000  0.350000  7.850000 0.680000 ;
      RECT  7.510000  1.745000  7.850000 1.765000 ;
      RECT  7.510000  1.765000  7.680000 2.375000 ;
      RECT  7.640000  0.680000  7.850000 1.575000 ;
      RECT  7.950000  1.915000  8.280000 2.425000 ;
      RECT  8.030000  0.345000  8.280000 1.055000 ;
      RECT  8.030000  1.055000 10.555000 1.275000 ;
      RECT  8.030000  1.275000  8.280000 1.915000 ;
      RECT  8.460000  0.085000  8.745000 0.545000 ;
      RECT  8.460000  1.835000  8.745000 2.635000 ;
      RECT  9.340000  0.085000  9.595000 0.545000 ;
      RECT  9.340000  1.810000  9.595000 2.635000 ;
      RECT 10.105000  0.085000 10.435000 0.545000 ;
      RECT 10.105000  1.810000 10.435000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.615000  1.785000  0.785000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  0.765000  1.235000 0.935000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.785000  2.615000 1.955000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  0.765000  3.075000 0.935000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.225000  1.105000  5.395000 1.275000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.555000 1.755000 0.845000 1.800000 ;
      RECT 0.555000 1.800000 5.435000 1.940000 ;
      RECT 0.555000 1.940000 0.845000 1.985000 ;
      RECT 1.005000 0.735000 1.295000 0.780000 ;
      RECT 1.005000 0.780000 3.135000 0.920000 ;
      RECT 1.005000 0.920000 1.295000 0.965000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.845000 0.735000 3.135000 0.780000 ;
      RECT 2.845000 0.920000 3.135000 0.965000 ;
      RECT 2.920000 0.965000 3.135000 1.120000 ;
      RECT 2.920000 1.120000 5.455000 1.260000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 5.165000 1.075000 5.455000 1.120000 ;
      RECT 5.165000 1.260000 5.455000 1.305000 ;
  END
END sky130_fd_sc_hd__dfstp_4
MACRO sky130_fd_sc_hd__dfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.005000 2.180000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.945000 0.265000 9.200000 0.795000 ;
        RECT 8.945000 1.655000 9.200000 2.325000 ;
        RECT 9.020000 0.795000 9.200000 1.655000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 0.735000 4.020000 1.065000 ;
      LAYER mcon ;
        RECT 3.850000 0.765000 4.020000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.680000 0.735000 7.340000 1.005000 ;
        RECT 6.680000 1.005000 7.010000 1.065000 ;
      LAYER mcon ;
        RECT 7.110000 0.765000 7.280000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.790000 0.735000 4.080000 0.780000 ;
        RECT 3.790000 0.780000 7.340000 0.920000 ;
        RECT 3.790000 0.920000 4.080000 0.965000 ;
        RECT 7.050000 0.735000 7.340000 0.780000 ;
        RECT 7.050000 0.920000 7.340000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.240000 2.465000 ;
      RECT 1.430000  0.635000 2.125000 0.825000 ;
      RECT 1.430000  0.825000 1.600000 1.795000 ;
      RECT 1.430000  1.795000 2.125000 1.965000 ;
      RECT 1.455000  0.085000 1.785000 0.465000 ;
      RECT 1.455000  2.135000 1.785000 2.635000 ;
      RECT 1.955000  0.305000 2.125000 0.635000 ;
      RECT 1.955000  1.965000 2.125000 2.465000 ;
      RECT 2.350000  0.705000 2.570000 1.575000 ;
      RECT 2.350000  1.575000 2.850000 1.955000 ;
      RECT 2.360000  2.250000 3.190000 2.420000 ;
      RECT 2.425000  0.265000 3.440000 0.465000 ;
      RECT 2.750000  0.645000 3.100000 1.015000 ;
      RECT 3.020000  1.195000 3.440000 1.235000 ;
      RECT 3.020000  1.235000 4.370000 1.405000 ;
      RECT 3.020000  1.405000 3.190000 2.250000 ;
      RECT 3.270000  0.465000 3.440000 1.195000 ;
      RECT 3.360000  1.575000 3.610000 1.835000 ;
      RECT 3.360000  1.835000 4.730000 2.085000 ;
      RECT 3.430000  2.255000 3.810000 2.635000 ;
      RECT 3.610000  0.085000 4.020000 0.525000 ;
      RECT 3.990000  2.085000 4.160000 2.375000 ;
      RECT 4.120000  1.405000 4.370000 1.565000 ;
      RECT 4.310000  0.295000 4.560000 0.725000 ;
      RECT 4.310000  0.725000 4.730000 1.065000 ;
      RECT 4.330000  2.255000 4.660000 2.635000 ;
      RECT 4.540000  1.065000 4.730000 1.835000 ;
      RECT 4.760000  0.085000 5.080000 0.545000 ;
      RECT 4.900000  0.725000 6.150000 0.895000 ;
      RECT 4.900000  0.895000 5.070000 1.655000 ;
      RECT 4.900000  1.655000 5.420000 1.965000 ;
      RECT 5.130000  2.165000 5.760000 2.415000 ;
      RECT 5.240000  1.065000 5.420000 1.475000 ;
      RECT 5.590000  1.235000 7.490000 1.405000 ;
      RECT 5.590000  1.405000 5.760000 1.915000 ;
      RECT 5.590000  1.915000 6.800000 2.085000 ;
      RECT 5.590000  2.085000 5.760000 2.165000 ;
      RECT 5.640000  0.305000 6.490000 0.475000 ;
      RECT 5.820000  0.895000 6.150000 1.015000 ;
      RECT 5.930000  1.575000 7.850000 1.745000 ;
      RECT 5.940000  2.255000 6.360000 2.635000 ;
      RECT 6.320000  0.475000 6.490000 1.235000 ;
      RECT 6.560000  2.085000 6.800000 2.375000 ;
      RECT 6.690000  0.085000 7.350000 0.565000 ;
      RECT 7.030000  1.945000 7.360000 2.635000 ;
      RECT 7.160000  1.175000 7.490000 1.235000 ;
      RECT 7.530000  0.350000 7.850000 0.680000 ;
      RECT 7.530000  1.745000 7.850000 1.765000 ;
      RECT 7.530000  1.765000 7.700000 2.375000 ;
      RECT 7.660000  0.680000 7.850000 1.575000 ;
      RECT 7.970000  1.915000 8.300000 2.425000 ;
      RECT 8.050000  0.345000 8.300000 0.995000 ;
      RECT 8.050000  0.995000 8.850000 1.325000 ;
      RECT 8.050000  1.325000 8.300000 1.915000 ;
      RECT 8.480000  0.085000 8.765000 0.545000 ;
      RECT 8.480000  1.835000 8.765000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.785000 0.780000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  0.765000 1.240000 0.935000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.785000 2.640000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  0.765000 3.100000 0.935000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.250000  1.105000 5.420000 1.275000 ;
      RECT 5.250000  1.785000 5.420000 1.955000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.755000 0.840000 1.800000 ;
      RECT 0.550000 1.800000 5.480000 1.940000 ;
      RECT 0.550000 1.940000 0.840000 1.985000 ;
      RECT 1.010000 0.735000 1.300000 0.780000 ;
      RECT 1.010000 0.780000 3.160000 0.920000 ;
      RECT 1.010000 0.920000 1.300000 0.965000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 0.735000 3.160000 0.780000 ;
      RECT 2.870000 0.920000 3.160000 0.965000 ;
      RECT 2.945000 0.965000 3.160000 1.120000 ;
      RECT 2.945000 1.120000 5.480000 1.260000 ;
      RECT 5.190000 1.075000 5.480000 1.120000 ;
      RECT 5.190000 1.260000 5.480000 1.305000 ;
      RECT 5.190000 1.755000 5.480000 1.800000 ;
      RECT 5.190000 1.940000 5.480000 1.985000 ;
  END
END sky130_fd_sc_hd__dfstp_1
MACRO sky130_fd_sc_hd__macro_sparecell
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__macro_sparecell ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.34000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN LO
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.215000 1.075000 4.965000 1.325000 ;
      LAYER mcon ;
        RECT 4.775000 1.105000 4.945000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.135000 1.075000 5.895000 1.325000 ;
      LAYER mcon ;
        RECT 5.705000 1.105000 5.875000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.755000 0.915000 7.275000 2.465000 ;
      LAYER mcon ;
        RECT 6.765000 1.105000 6.935000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.445000 1.075000 8.205000 1.325000 ;
      LAYER mcon ;
        RECT 7.625000 1.105000 7.795000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.375000 1.075000 9.125000 1.325000 ;
      LAYER mcon ;
        RECT 8.485000 1.105000 8.655000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.715000 1.075000 5.005000 1.120000 ;
        RECT 4.715000 1.120000 8.715000 1.260000 ;
        RECT 4.715000 1.260000 5.005000 1.305000 ;
        RECT 5.645000 1.075000 5.935000 1.120000 ;
        RECT 5.645000 1.260000 5.935000 1.305000 ;
        RECT 6.705000 1.075000 6.995000 1.120000 ;
        RECT 6.705000 1.260000 6.995000 1.305000 ;
        RECT 7.565000 1.075000 7.855000 1.120000 ;
        RECT 7.565000 1.260000 7.855000 1.305000 ;
        RECT 8.425000 1.075000 8.715000 1.120000 ;
        RECT 8.425000 1.260000 8.715000 1.305000 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.340000 0.085000 ;
        RECT  0.145000  0.085000  0.355000 0.905000 ;
        RECT  1.025000  0.085000  1.255000 0.905000 ;
        RECT  1.515000  0.085000  1.805000 0.555000 ;
        RECT  2.475000  0.085000  2.645000 0.555000 ;
        RECT  3.315000  0.085000  3.590000 0.905000 ;
        RECT  5.215000  0.085000  5.385000 0.545000 ;
        RECT  6.755000  0.085000  7.095000 0.745000 ;
        RECT  7.955000  0.085000  8.125000 0.545000 ;
        RECT  9.750000  0.085000 10.025000 0.905000 ;
        RECT 10.695000  0.085000 10.865000 0.555000 ;
        RECT 11.535000  0.085000 11.825000 0.555000 ;
        RECT 12.085000  0.085000 12.315000 0.905000 ;
        RECT 12.985000  0.085000 13.195000 0.905000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
        RECT 11.645000 -0.085000 11.815000 0.085000 ;
        RECT 12.105000 -0.085000 12.275000 0.085000 ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
        RECT 13.025000 -0.085000 13.195000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 13.530000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 13.340000 2.805000 ;
        RECT  0.145000 1.495000  0.355000 2.635000 ;
        RECT  1.025000 1.495000  1.255000 2.635000 ;
        RECT  2.815000 1.835000  3.145000 2.635000 ;
        RECT  3.870000 1.835000  4.125000 2.635000 ;
        RECT  4.795000 1.835000  4.965000 2.635000 ;
        RECT  5.635000 1.495000  5.895000 2.635000 ;
        RECT  6.255000 1.910000  6.585000 2.635000 ;
        RECT  7.445000 1.495000  7.705000 2.635000 ;
        RECT  8.375000 1.835000  8.545000 2.635000 ;
        RECT  9.215000 1.835000  9.470000 2.635000 ;
        RECT 10.195000 1.835000 10.525000 2.635000 ;
        RECT 12.085000 1.495000 12.315000 2.635000 ;
        RECT 12.985000 1.495000 13.195000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
        RECT 11.185000 2.635000 11.355000 2.805000 ;
        RECT 11.645000 2.635000 11.815000 2.805000 ;
        RECT 12.105000 2.635000 12.275000 2.805000 ;
        RECT 12.565000 2.635000 12.735000 2.805000 ;
        RECT 13.025000 2.635000 13.195000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.525000 0.255000  0.855000 0.885000 ;
      RECT  0.525000 0.885000  0.775000 1.485000 ;
      RECT  0.525000 1.485000  0.855000 2.465000 ;
      RECT  0.945000 1.075000  1.275000 1.325000 ;
      RECT  1.505000 1.835000  1.805000 2.295000 ;
      RECT  1.505000 2.295000  2.645000 2.465000 ;
      RECT  1.545000 0.735000  3.145000 0.905000 ;
      RECT  1.545000 0.905000  1.760000 1.445000 ;
      RECT  1.545000 1.445000  2.305000 1.665000 ;
      RECT  1.930000 1.075000  2.700000 1.275000 ;
      RECT  1.975000 0.255000  2.305000 0.725000 ;
      RECT  1.975000 0.725000  3.145000 0.735000 ;
      RECT  1.975000 1.665000  2.305000 2.125000 ;
      RECT  2.475000 1.455000  3.590000 1.665000 ;
      RECT  2.475000 1.665000  2.645000 2.295000 ;
      RECT  2.815000 0.255000  3.145000 0.725000 ;
      RECT  2.870000 1.075000  3.590000 1.275000 ;
      RECT  3.315000 1.665000  3.590000 2.465000 ;
      RECT  3.765000 0.655000  4.625000 0.905000 ;
      RECT  3.765000 0.905000  4.045000 1.495000 ;
      RECT  3.765000 1.495000  5.465000 1.665000 ;
      RECT  3.875000 0.255000  5.045000 0.465000 ;
      RECT  3.875000 0.465000  4.205000 0.485000 ;
      RECT  4.295000 1.665000  4.625000 2.465000 ;
      RECT  4.795000 0.465000  5.045000 0.715000 ;
      RECT  4.795000 0.715000  5.895000 0.885000 ;
      RECT  5.135000 1.665000  5.465000 2.465000 ;
      RECT  5.555000 0.255000  5.895000 0.715000 ;
      RECT  6.065000 0.255000  6.585000 1.740000 ;
      RECT  7.445000 0.255000  7.785000 0.715000 ;
      RECT  7.445000 0.715000  8.545000 0.885000 ;
      RECT  7.875000 1.495000  9.575000 1.665000 ;
      RECT  7.875000 1.665000  8.205000 2.465000 ;
      RECT  8.295000 0.255000  9.465000 0.465000 ;
      RECT  8.295000 0.465000  8.545000 0.715000 ;
      RECT  8.715000 0.655000  9.575000 0.905000 ;
      RECT  8.715000 1.665000  9.045000 2.465000 ;
      RECT  9.135000 0.465000  9.465000 0.485000 ;
      RECT  9.295000 0.905000  9.575000 1.495000 ;
      RECT  9.750000 1.075000 10.470000 1.275000 ;
      RECT  9.750000 1.455000 10.865000 1.665000 ;
      RECT  9.750000 1.665000 10.025000 2.465000 ;
      RECT 10.195000 0.255000 10.525000 0.725000 ;
      RECT 10.195000 0.725000 11.365000 0.735000 ;
      RECT 10.195000 0.735000 11.795000 0.905000 ;
      RECT 10.640000 1.075000 11.410000 1.275000 ;
      RECT 10.695000 1.665000 10.865000 2.295000 ;
      RECT 10.695000 2.295000 11.835000 2.465000 ;
      RECT 11.035000 0.255000 11.365000 0.725000 ;
      RECT 11.035000 1.445000 11.795000 1.665000 ;
      RECT 11.035000 1.665000 11.365000 2.125000 ;
      RECT 11.535000 1.835000 11.835000 2.295000 ;
      RECT 11.580000 0.905000 11.795000 1.445000 ;
      RECT 12.065000 1.075000 12.395000 1.325000 ;
      RECT 12.485000 0.255000 12.815000 0.885000 ;
      RECT 12.485000 1.485000 12.815000 2.465000 ;
      RECT 12.565000 0.885000 12.815000 1.485000 ;
    LAYER mcon ;
      RECT  0.565000 1.105000  0.735000 1.275000 ;
      RECT  1.085000 1.105000  1.255000 1.275000 ;
      RECT  1.570000 1.105000  1.740000 1.275000 ;
      RECT  2.100000 1.105000  2.270000 1.275000 ;
      RECT  2.960000 1.105000  3.130000 1.275000 ;
      RECT  3.820000 1.105000  3.990000 1.275000 ;
      RECT  9.345000 1.105000  9.515000 1.275000 ;
      RECT 10.205000 1.105000 10.375000 1.275000 ;
      RECT 11.065000 1.105000 11.235000 1.275000 ;
      RECT 11.605000 1.105000 11.775000 1.275000 ;
      RECT 12.090000 1.105000 12.260000 1.275000 ;
      RECT 12.605000 1.105000 12.775000 1.275000 ;
    LAYER met1 ;
      RECT  0.505000 1.075000  0.875000 1.305000 ;
      RECT  1.025000 1.075000  1.315000 1.120000 ;
      RECT  1.025000 1.120000  1.800000 1.260000 ;
      RECT  1.025000 1.260000  1.315000 1.305000 ;
      RECT  1.510000 1.075000  1.800000 1.120000 ;
      RECT  1.510000 1.260000  1.800000 1.305000 ;
      RECT  2.040000 1.075000  2.330000 1.120000 ;
      RECT  2.040000 1.120000  4.050000 1.260000 ;
      RECT  2.040000 1.260000  2.330000 1.305000 ;
      RECT  2.900000 1.075000  3.190000 1.120000 ;
      RECT  2.900000 1.260000  3.190000 1.305000 ;
      RECT  3.760000 1.075000  4.050000 1.120000 ;
      RECT  3.760000 1.260000  4.050000 1.305000 ;
      RECT  9.285000 1.075000  9.575000 1.120000 ;
      RECT  9.285000 1.120000 11.295000 1.260000 ;
      RECT  9.285000 1.260000  9.575000 1.305000 ;
      RECT 10.145000 1.075000 10.435000 1.120000 ;
      RECT 10.145000 1.260000 10.435000 1.305000 ;
      RECT 11.005000 1.075000 11.295000 1.120000 ;
      RECT 11.005000 1.260000 11.295000 1.305000 ;
      RECT 11.545000 1.075000 11.835000 1.120000 ;
      RECT 11.545000 1.120000 12.320000 1.260000 ;
      RECT 11.545000 1.260000 11.835000 1.305000 ;
      RECT 12.030000 1.075000 12.320000 1.120000 ;
      RECT 12.030000 1.260000 12.320000 1.305000 ;
      RECT 12.470000 1.075000 12.835000 1.305000 ;
    LAYER pwell ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  3.360000 -0.085000  3.530000 0.085000 ;
      RECT  5.660000 -0.085000  5.830000 0.085000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  7.510000 -0.085000  7.680000 0.085000 ;
      RECT  9.810000 -0.085000  9.980000 0.085000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
  END
END sky130_fd_sc_hd__macro_sparecell
MACRO sky130_fd_sc_hd__lpflow_isobufsrckapwr_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.26000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.615000 1.320000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.260000 1.075000 4.700000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.340000 0.280000  7.600000 0.735000 ;
        RECT  7.340000 0.735000 14.085000 0.905000 ;
        RECT  7.375000 1.495000 14.085000 1.720000 ;
        RECT  7.375000 1.720000 12.745000 1.735000 ;
        RECT  7.375000 1.735000  7.600000 2.460000 ;
        RECT  8.200000 0.280000  8.460000 0.735000 ;
        RECT  8.200000 1.735000  8.460000 2.460000 ;
        RECT  9.060000 0.280000  9.320000 0.735000 ;
        RECT  9.060000 1.735000  9.320000 2.460000 ;
        RECT  9.905000 0.280000 10.180000 0.735000 ;
        RECT  9.920000 1.735000 10.180000 2.460000 ;
        RECT 10.765000 0.280000 11.025000 0.735000 ;
        RECT 10.765000 1.735000 11.025000 2.460000 ;
        RECT 11.625000 0.280000 11.885000 0.735000 ;
        RECT 11.625000 1.735000 11.885000 2.460000 ;
        RECT 12.485000 0.280000 12.745000 0.735000 ;
        RECT 12.485000 1.735000 12.745000 2.460000 ;
        RECT 12.920000 0.905000 14.085000 1.495000 ;
        RECT 13.355000 0.280000 13.615000 0.735000 ;
        RECT 13.355000 1.720000 13.645000 2.460000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 10.350000 1.905000 10.595000 2.465000 ;
      LAYER mcon ;
        RECT 10.395000 2.125000 10.565000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 11.210000 1.905000 11.455000 2.465000 ;
      LAYER mcon ;
        RECT 11.255000 2.125000 11.425000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 12.070000 1.905000 12.315000 2.465000 ;
      LAYER mcon ;
        RECT 12.110000 2.125000 12.280000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 12.930000 1.905000 13.185000 2.465000 ;
      LAYER mcon ;
        RECT 12.960000 2.125000 13.130000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 13.815000 1.890000 14.085000 2.465000 ;
      LAYER mcon ;
        RECT 13.840000 2.125000 14.010000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.155000 1.495000 5.485000 2.465000 ;
      LAYER mcon ;
        RECT 5.235000 2.125000 5.405000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.015000 1.495000 6.345000 2.465000 ;
      LAYER mcon ;
        RECT 6.095000 2.125000 6.265000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.875000 1.495000 7.205000 2.465000 ;
      LAYER mcon ;
        RECT 6.950000 2.125000 7.120000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.770000 1.905000 8.030000 2.465000 ;
      LAYER mcon ;
        RECT 7.800000 2.125000 7.970000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.630000 1.905000 8.890000 2.465000 ;
      LAYER mcon ;
        RECT 8.680000 2.125000 8.850000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.490000 1.905000 9.750000 2.465000 ;
      LAYER mcon ;
        RECT 9.540000 2.125000 9.710000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT  0.070000 2.140000 14.190000 2.340000 ;
        RECT  5.175000 2.080000  5.465000 2.140000 ;
        RECT  6.035000 2.080000  6.325000 2.140000 ;
        RECT  6.890000 2.080000  7.180000 2.140000 ;
        RECT  7.740000 2.080000  8.030000 2.140000 ;
        RECT  8.620000 2.080000  8.910000 2.140000 ;
        RECT  9.480000 2.080000  9.770000 2.140000 ;
        RECT 10.335000 2.080000 10.625000 2.140000 ;
        RECT 11.195000 2.080000 11.485000 2.140000 ;
        RECT 12.050000 2.080000 12.340000 2.140000 ;
        RECT 12.900000 2.080000 13.190000 2.140000 ;
        RECT 13.780000 2.080000 14.070000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
    PORT
      LAYER pwell ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 14.450000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.130000  1.495000  0.535000 2.635000 ;
      RECT  0.245000  0.085000  0.535000 0.905000 ;
      RECT  0.705000  0.255000  1.035000 0.815000 ;
      RECT  0.705000  1.575000  1.035000 2.465000 ;
      RECT  0.785000  0.815000  1.035000 1.075000 ;
      RECT  0.785000  1.075000  2.265000 1.275000 ;
      RECT  0.785000  1.275000  1.035000 1.575000 ;
      RECT  1.205000  1.575000  1.585000 2.295000 ;
      RECT  1.205000  2.295000  3.265000 2.465000 ;
      RECT  1.215000  0.085000  1.505000 0.905000 ;
      RECT  1.675000  0.255000  2.005000 0.725000 ;
      RECT  1.675000  0.725000  4.525000 0.905000 ;
      RECT  1.755000  1.445000  2.765000 1.745000 ;
      RECT  1.755000  1.745000  1.925000 2.125000 ;
      RECT  2.095000  1.935000  2.425000 2.295000 ;
      RECT  2.175000  0.085000  2.345000 0.555000 ;
      RECT  2.435000  0.905000  3.095000 0.965000 ;
      RECT  2.435000  0.965000  2.765000 1.445000 ;
      RECT  2.515000  0.255000  2.845000 0.725000 ;
      RECT  2.595000  1.745000  2.765000 2.125000 ;
      RECT  2.935000  1.455000  4.975000 1.665000 ;
      RECT  2.935000  1.665000  3.265000 2.295000 ;
      RECT  3.015000  0.085000  3.185000 0.555000 ;
      RECT  3.355000  0.255000  3.685000 0.725000 ;
      RECT  3.435000  1.835000  3.685000 2.635000 ;
      RECT  3.855000  0.085000  4.025000 0.555000 ;
      RECT  3.855000  1.665000  4.025000 2.465000 ;
      RECT  4.195000  0.255000  4.525000 0.725000 ;
      RECT  4.195000  1.835000  4.525000 2.635000 ;
      RECT  4.695000  0.085000  5.450000 0.565000 ;
      RECT  4.695000  0.565000  4.975000 0.905000 ;
      RECT  4.695000  1.665000  4.975000 2.465000 ;
      RECT  5.145000  0.735000  5.460000 1.325000 ;
      RECT  5.655000  0.265000  5.880000 1.075000 ;
      RECT  5.655000  1.075000 12.750000 1.325000 ;
      RECT  5.655000  1.325000  5.845000 2.465000 ;
      RECT  6.050000  0.085000  6.310000 0.610000 ;
      RECT  6.490000  0.265000  6.740000 1.075000 ;
      RECT  6.515000  1.325000  6.705000 2.460000 ;
      RECT  6.910000  0.085000  7.170000 0.645000 ;
      RECT  7.770000  0.085000  8.030000 0.565000 ;
      RECT  8.630000  0.085000  8.890000 0.565000 ;
      RECT  9.490000  0.085000  9.735000 0.565000 ;
      RECT 10.350000  0.085000 10.595000 0.565000 ;
      RECT 11.205000  0.085000 11.455000 0.565000 ;
      RECT 12.065000  0.085000 12.315000 0.565000 ;
      RECT 12.925000  0.085000 13.185000 0.565000 ;
      RECT 13.785000  0.085000 14.085000 0.565000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.525000  0.765000  2.695000 0.935000 ;
      RECT  2.885000  0.765000  3.055000 0.935000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.210000  0.765000  5.380000 0.935000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT 2.465000 0.735000 3.115000 0.780000 ;
      RECT 2.465000 0.780000 5.440000 0.920000 ;
      RECT 2.465000 0.920000 3.115000 0.965000 ;
      RECT 5.150000 0.735000 5.440000 0.780000 ;
      RECT 5.150000 0.920000 5.440000 0.965000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrckapwr_16
MACRO sky130_fd_sc_hd__mux2i_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2i_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.060000 0.420000 1.285000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 0.995000 1.125000 1.155000 ;
        RECT 0.955000 1.155000 1.205000 1.325000 ;
        RECT 1.035000 1.325000 1.205000 1.445000 ;
        RECT 1.035000 1.445000 1.235000 2.110000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.260000 0.760000 3.595000 1.620000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 0.595000 0.780000 1.455000 ;
        RECT 0.590000 1.455000 0.840000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.255000 1.805000 0.425000 ;
      RECT 0.085000  0.425000 0.440000 0.465000 ;
      RECT 0.085000  0.465000 0.345000 0.885000 ;
      RECT 0.120000  1.455000 0.420000 2.295000 ;
      RECT 0.120000  2.295000 1.575000 2.465000 ;
      RECT 0.955000  0.655000 1.520000 0.715000 ;
      RECT 0.955000  0.715000 2.620000 0.825000 ;
      RECT 0.965000  0.425000 1.805000 0.465000 ;
      RECT 1.295000  0.825000 2.620000 0.885000 ;
      RECT 1.385000  1.075000 3.085000 1.310000 ;
      RECT 1.405000  1.480000 2.615000 1.650000 ;
      RECT 1.405000  1.650000 1.575000 2.295000 ;
      RECT 1.745000  1.835000 1.975000 2.635000 ;
      RECT 1.975000  0.085000 2.145000 0.545000 ;
      RECT 2.285000  1.650000 2.615000 2.465000 ;
      RECT 2.385000  0.255000 2.620000 0.715000 ;
      RECT 2.800000  0.255000 3.165000 0.485000 ;
      RECT 2.800000  0.485000 3.085000 1.075000 ;
      RECT 2.860000  1.310000 3.085000 2.465000 ;
      RECT 3.295000  1.835000 3.590000 2.635000 ;
      RECT 3.335000  0.085000 3.555000 0.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__mux2i_1
MACRO sky130_fd_sc_hd__mux2i_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2i_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 1.075000 3.560000 1.275000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.310000 0.995000 4.635000 1.615000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.780000 1.325000 ;
        RECT 0.580000 0.725000 0.780000 0.995000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  1.691250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715000 0.295000 4.975000 0.465000 ;
        RECT 2.715000 2.255000 4.975000 2.425000 ;
        RECT 4.750000 1.785000 4.975000 2.255000 ;
        RECT 4.805000 0.465000 4.975000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.675000 ;
      RECT 0.085000  0.675000 0.260000 1.495000 ;
      RECT 0.085000  1.495000 1.395000 1.665000 ;
      RECT 0.085000  1.665000 0.260000 2.135000 ;
      RECT 0.085000  2.135000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.835000 0.545000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 0.935000  1.835000 1.735000 2.005000 ;
      RECT 1.015000  0.575000 1.255000 0.935000 ;
      RECT 1.225000  1.155000 1.985000 1.325000 ;
      RECT 1.225000  1.325000 1.395000 1.495000 ;
      RECT 1.355000  2.255000 1.685000 2.635000 ;
      RECT 1.435000  0.085000 1.685000 0.885000 ;
      RECT 1.565000  1.495000 3.465000 1.665000 ;
      RECT 1.565000  1.665000 1.735000 1.835000 ;
      RECT 1.655000  1.075000 1.985000 1.155000 ;
      RECT 1.855000  0.295000 2.025000 0.735000 ;
      RECT 1.855000  0.735000 3.465000 0.905000 ;
      RECT 1.855000  2.135000 2.080000 2.465000 ;
      RECT 1.910000  1.835000 2.885000 1.915000 ;
      RECT 1.910000  1.915000 4.350000 2.005000 ;
      RECT 1.910000  2.005000 2.080000 2.135000 ;
      RECT 2.275000  0.085000 2.445000 0.545000 ;
      RECT 2.275000  2.175000 2.525000 2.635000 ;
      RECT 2.715000  2.005000 4.350000 2.085000 ;
      RECT 3.135000  0.655000 3.465000 0.735000 ;
      RECT 3.135000  1.665000 3.465000 1.715000 ;
      RECT 3.850000  0.655000 4.345000 0.825000 ;
      RECT 3.850000  0.825000 4.105000 0.935000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  0.765000 1.240000 0.935000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 3.850000  0.765000 4.020000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
    LAYER met1 ;
      RECT 1.010000 0.735000 1.300000 0.780000 ;
      RECT 1.010000 0.780000 4.080000 0.920000 ;
      RECT 1.010000 0.920000 1.300000 0.965000 ;
      RECT 3.790000 0.735000 4.080000 0.780000 ;
      RECT 3.790000 0.920000 4.080000 0.965000 ;
  END
END sky130_fd_sc_hd__mux2i_2
MACRO sky130_fd_sc_hd__mux2i_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2i_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 0.995000 1.070000 1.105000 ;
        RECT 0.560000 1.105000 1.240000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 0.995000 3.550000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.237500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.845000 1.075000 5.930000 1.290000 ;
        RECT 5.760000 1.290000 5.930000 1.425000 ;
        RECT 5.760000 1.425000 7.850000 1.595000 ;
        RECT 7.680000 0.995000 7.850000 1.425000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  2.194500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.315000 3.785000 0.485000 ;
        RECT 0.095000 0.485000 0.320000 2.255000 ;
        RECT 0.095000 2.255000 3.785000 2.425000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.515000  0.655000 1.700000 0.825000 ;
      RECT 0.515000  1.575000 5.580000 1.745000 ;
      RECT 1.355000  0.825000 1.700000 0.935000 ;
      RECT 2.195000  0.655000 5.485000 0.825000 ;
      RECT 2.195000  1.915000 7.165000 2.085000 ;
      RECT 3.975000  0.085000 4.305000 0.465000 ;
      RECT 3.975000  2.255000 4.305000 2.635000 ;
      RECT 4.475000  0.255000 4.645000 0.655000 ;
      RECT 4.815000  0.085000 5.145000 0.465000 ;
      RECT 4.815000  2.255000 5.145000 2.635000 ;
      RECT 5.315000  0.255000 5.485000 0.655000 ;
      RECT 5.655000  0.085000 5.980000 0.590000 ;
      RECT 5.655000  2.255000 5.985000 2.635000 ;
      RECT 6.150000  0.255000 6.325000 0.715000 ;
      RECT 6.150000  0.715000 7.165000 0.905000 ;
      RECT 6.150000  0.905000 6.450000 0.935000 ;
      RECT 6.155000  1.795000 6.325000 1.915000 ;
      RECT 6.155000  2.085000 6.325000 2.465000 ;
      RECT 6.495000  2.255000 6.825000 2.635000 ;
      RECT 6.545000  0.085000 6.795000 0.545000 ;
      RECT 6.730000  1.075000 7.510000 1.245000 ;
      RECT 6.995000  0.510000 7.165000 0.715000 ;
      RECT 6.995000  1.795000 7.165000 1.915000 ;
      RECT 6.995000  2.085000 7.165000 2.465000 ;
      RECT 7.340000  0.655000 8.195000 0.825000 ;
      RECT 7.340000  0.825000 7.510000 1.075000 ;
      RECT 7.435000  0.085000 7.765000 0.465000 ;
      RECT 7.435000  2.255000 7.765000 2.635000 ;
      RECT 7.935000  0.255000 8.195000 0.655000 ;
      RECT 7.935000  1.795000 8.195000 2.465000 ;
      RECT 8.020000  0.825000 8.195000 1.795000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.530000  0.765000 1.700000 0.935000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.150000  0.765000 6.320000 0.935000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 1.470000 0.735000 1.760000 0.780000 ;
      RECT 1.470000 0.780000 6.380000 0.920000 ;
      RECT 1.470000 0.920000 1.760000 0.965000 ;
      RECT 6.090000 0.735000 6.380000 0.780000 ;
      RECT 6.090000 0.920000 6.380000 0.965000 ;
  END
END sky130_fd_sc_hd__mux2i_4
MACRO sky130_fd_sc_hd__fah_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fah_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.42000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 1.075000 1.440000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.691500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.075000 2.495000 1.275000 ;
        RECT 1.990000 1.275000 2.190000 1.410000 ;
        RECT 2.015000 1.410000 2.190000 1.725000 ;
      LAYER mcon ;
        RECT 1.990000 1.105000 2.160000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.675000 0.995000 5.925000 1.325000 ;
      LAYER mcon ;
        RECT 5.680000 1.105000 5.850000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.930000 1.075000 2.220000 1.120000 ;
        RECT 1.930000 1.120000 5.910000 1.260000 ;
        RECT 1.930000 1.260000 2.220000 1.305000 ;
        RECT 5.620000 1.075000 5.910000 1.120000 ;
        RECT 5.620000 1.260000 5.910000 1.305000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.475000 1.075000  9.865000 1.325000 ;
        RECT 9.690000 0.735000 10.010000 0.935000 ;
        RECT 9.690000 0.935000  9.865000 1.075000 ;
    END
  END CI
  PIN COUT
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.870000 0.270000 11.310000 0.825000 ;
        RECT 10.870000 0.825000 11.040000 1.495000 ;
        RECT 10.870000 1.495000 11.390000 2.465000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.506000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.980000 0.255000 12.335000 0.825000 ;
        RECT 11.985000 1.785000 12.335000 2.465000 ;
        RECT 12.110000 0.825000 12.335000 1.785000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.610000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.085000  0.255000  0.425000 0.805000 ;
      RECT  0.085000  0.805000  0.255000 1.500000 ;
      RECT  0.085000  1.500000  0.445000 1.895000 ;
      RECT  0.085000  1.895000  2.805000 2.065000 ;
      RECT  0.085000  2.065000  0.395000 2.465000 ;
      RECT  0.425000  0.995000  0.780000 1.325000 ;
      RECT  0.565000  2.260000  0.930000 2.635000 ;
      RECT  0.595000  0.085000  0.765000 0.545000 ;
      RECT  0.595000  0.735000  1.320000 0.905000 ;
      RECT  0.595000  0.905000  0.780000 0.995000 ;
      RECT  0.610000  1.325000  0.780000 1.380000 ;
      RECT  0.610000  1.380000  0.815000 1.445000 ;
      RECT  0.610000  1.445000  1.315000 1.455000 ;
      RECT  0.615000  1.455000  1.315000 1.615000 ;
      RECT  0.985000  1.615000  1.315000 1.715000 ;
      RECT  0.990000  0.255000  1.320000 0.735000 ;
      RECT  1.490000  1.445000  1.820000 1.500000 ;
      RECT  1.490000  1.500000  1.840000 1.725000 ;
      RECT  1.500000  0.255000  1.840000 0.715000 ;
      RECT  1.500000  0.715000  2.520000 0.885000 ;
      RECT  1.500000  0.885000  1.820000 0.905000 ;
      RECT  1.615000  0.905000  1.820000 1.445000 ;
      RECT  2.010000  0.085000  2.180000 0.545000 ;
      RECT  2.065000  2.235000  2.395000 2.635000 ;
      RECT  2.350000  0.255000  4.840000 0.425000 ;
      RECT  2.350000  0.425000  2.520000 0.715000 ;
      RECT  2.360000  1.445000  2.860000 1.715000 ;
      RECT  2.635000  2.065000  2.805000 2.295000 ;
      RECT  2.635000  2.295000  4.950000 2.465000 ;
      RECT  2.690000  0.595000  2.860000 1.445000 ;
      RECT  3.030000  0.425000  4.840000 0.465000 ;
      RECT  3.030000  0.465000  3.200000 1.955000 ;
      RECT  3.030000  1.955000  4.320000 2.125000 ;
      RECT  3.370000  0.635000  3.900000 0.805000 ;
      RECT  3.370000  0.805000  3.540000 1.455000 ;
      RECT  3.370000  1.455000  3.815000 1.785000 ;
      RECT  3.985000  1.785000  4.320000 1.955000 ;
      RECT  4.070000  0.645000  4.400000 0.735000 ;
      RECT  4.070000  0.735000  4.560000 0.755000 ;
      RECT  4.070000  0.755000  5.170000 0.780000 ;
      RECT  4.070000  0.780000  5.155000 0.805000 ;
      RECT  4.070000  0.805000  5.145000 0.905000 ;
      RECT  4.070000  1.075000  4.400000 1.160000 ;
      RECT  4.070000  1.160000  4.535000 1.615000 ;
      RECT  4.480000  0.905000  5.145000 0.925000 ;
      RECT  4.650000  0.465000  4.840000 0.585000 ;
      RECT  4.705000  0.925000  4.875000 2.295000 ;
      RECT  4.925000  0.735000  5.180000 0.740000 ;
      RECT  4.925000  0.740000  5.170000 0.755000 ;
      RECT  4.950000  0.715000  5.180000 0.735000 ;
      RECT  4.980000  0.690000  5.180000 0.715000 ;
      RECT  5.000000  0.655000  5.180000 0.690000 ;
      RECT  5.010000  0.255000  6.100000 0.425000 ;
      RECT  5.010000  0.425000  5.180000 0.655000 ;
      RECT  5.125000  1.150000  5.505000 1.320000 ;
      RECT  5.125000  1.320000  5.295000 2.295000 ;
      RECT  5.125000  2.295000  7.560000 2.465000 ;
      RECT  5.320000  0.865000  5.520000 0.925000 ;
      RECT  5.320000  0.925000  5.505000 1.150000 ;
      RECT  5.335000  0.840000  5.520000 0.865000 ;
      RECT  5.350000  0.595000  5.520000 0.840000 ;
      RECT  5.475000  1.700000  5.875000 2.030000 ;
      RECT  5.750000  0.425000  6.100000 0.565000 ;
      RECT  6.105000  0.740000  6.435000 1.275000 ;
      RECT  6.105000  1.445000  6.460000 1.615000 ;
      RECT  6.270000  0.255000  9.735000 0.425000 ;
      RECT  6.270000  0.425000  6.600000 0.570000 ;
      RECT  6.290000  1.615000  6.460000 1.955000 ;
      RECT  6.290000  1.955000  7.220000 2.125000 ;
      RECT  6.610000  0.755000  6.940000 0.925000 ;
      RECT  6.610000  0.925000  6.880000 1.275000 ;
      RECT  6.710000  1.275000  6.880000 1.785000 ;
      RECT  6.770000  0.595000  6.940000 0.755000 ;
      RECT  7.050000  1.060000  7.280000 1.130000 ;
      RECT  7.050000  1.130000  7.245000 1.175000 ;
      RECT  7.050000  1.175000  7.220000 1.955000 ;
      RECT  7.065000  1.045000  7.280000 1.060000 ;
      RECT  7.090000  1.010000  7.280000 1.045000 ;
      RECT  7.110000  0.595000  7.445000 0.765000 ;
      RECT  7.110000  0.765000  7.280000 1.010000 ;
      RECT  7.390000  1.275000  7.620000 1.375000 ;
      RECT  7.390000  1.375000  7.595000 1.400000 ;
      RECT  7.390000  1.400000  7.575000 1.425000 ;
      RECT  7.390000  1.425000  7.560000 2.295000 ;
      RECT  7.450000  0.995000  7.620000 1.275000 ;
      RECT  7.705000  0.425000  7.960000 0.825000 ;
      RECT  7.730000  1.510000  7.960000 2.295000 ;
      RECT  7.730000  2.295000  9.655000 2.465000 ;
      RECT  7.790000  0.825000  7.960000 1.510000 ;
      RECT  8.145000  1.955000  9.250000 2.125000 ;
      RECT  8.155000  0.595000  8.405000 0.925000 ;
      RECT  8.225000  0.925000  8.405000 1.445000 ;
      RECT  8.225000  1.445000  8.910000 1.785000 ;
      RECT  8.575000  0.595000  8.745000 1.105000 ;
      RECT  8.575000  1.105000  9.250000 1.275000 ;
      RECT  8.920000  0.685000  9.300000 0.935000 ;
      RECT  9.080000  1.275000  9.250000 1.955000 ;
      RECT  9.400000  0.425000  9.735000 0.515000 ;
      RECT  9.420000  1.495000 10.350000 1.705000 ;
      RECT  9.420000  1.705000  9.655000 2.295000 ;
      RECT  9.840000  2.275000 10.175000 2.635000 ;
      RECT  9.905000  0.085000 10.075000 0.565000 ;
      RECT 10.180000  0.995000 10.350000 1.495000 ;
      RECT 10.245000  0.285000 10.690000 0.825000 ;
      RECT 10.345000  1.875000 10.690000 2.465000 ;
      RECT 10.520000  0.825000 10.690000 1.875000 ;
      RECT 11.210000  0.995000 11.460000 1.325000 ;
      RECT 11.480000  0.085000 11.810000 0.825000 ;
      RECT 11.560000  1.785000 11.815000 2.635000 ;
      RECT 11.630000  0.995000 11.940000 1.615000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.450000  1.445000  2.620000 1.615000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.370000  0.765000  3.540000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.365000  1.445000  4.535000 1.615000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.570000  1.785000  5.740000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.150000  0.765000  6.320000 0.935000 ;
      RECT  6.150000  1.445000  6.320000 1.615000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.610000  1.105000  6.780000 1.275000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.460000  1.445000  8.630000 1.615000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.920000  0.765000  9.090000 0.935000 ;
      RECT  9.080000  1.785000  9.250000 1.955000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.520000  1.785000 10.690000 1.955000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.220000  1.105000 11.390000 1.275000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 11.680000  1.445000 11.850000 1.615000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
    LAYER met1 ;
      RECT  2.390000 1.415000  2.680000 1.460000 ;
      RECT  2.390000 1.460000  6.380000 1.600000 ;
      RECT  2.390000 1.600000  2.680000 1.645000 ;
      RECT  3.310000 0.735000  3.600000 0.780000 ;
      RECT  3.310000 0.780000  9.150000 0.920000 ;
      RECT  3.310000 0.920000  3.600000 0.965000 ;
      RECT  3.925000 1.755000  4.215000 1.800000 ;
      RECT  3.925000 1.800000  5.800000 1.940000 ;
      RECT  3.925000 1.940000  4.215000 1.985000 ;
      RECT  4.305000 1.415000  4.595000 1.460000 ;
      RECT  4.305000 1.600000  4.595000 1.645000 ;
      RECT  5.510000 1.755000  5.800000 1.800000 ;
      RECT  5.510000 1.940000  5.800000 1.985000 ;
      RECT  6.090000 0.735000  6.380000 0.780000 ;
      RECT  6.090000 0.920000  6.380000 0.965000 ;
      RECT  6.090000 1.415000  6.380000 1.460000 ;
      RECT  6.090000 1.600000  6.380000 1.645000 ;
      RECT  6.550000 1.075000  6.840000 1.120000 ;
      RECT  6.550000 1.120000 11.450000 1.260000 ;
      RECT  6.550000 1.260000  6.840000 1.305000 ;
      RECT  8.400000 1.415000  8.690000 1.460000 ;
      RECT  8.400000 1.460000 11.910000 1.600000 ;
      RECT  8.400000 1.600000  8.690000 1.645000 ;
      RECT  8.860000 0.735000  9.150000 0.780000 ;
      RECT  8.860000 0.920000  9.150000 0.965000 ;
      RECT  9.020000 1.755000  9.310000 1.800000 ;
      RECT  9.020000 1.800000 10.750000 1.940000 ;
      RECT  9.020000 1.940000  9.310000 1.985000 ;
      RECT 10.460000 1.755000 10.750000 1.800000 ;
      RECT 10.460000 1.940000 10.750000 1.985000 ;
      RECT 11.160000 1.075000 11.450000 1.120000 ;
      RECT 11.160000 1.260000 11.450000 1.305000 ;
      RECT 11.620000 1.415000 11.910000 1.460000 ;
      RECT 11.620000 1.600000 11.910000 1.645000 ;
  END
END sky130_fd_sc_hd__fah_1
MACRO sky130_fd_sc_hd__o2bb2a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.075000 3.645000 1.445000 ;
        RECT 3.315000 1.445000 4.965000 1.615000 ;
        RECT 4.605000 1.075000 4.965000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 1.075000 4.435000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.575000 1.445000 ;
        RECT 0.085000 1.445000 1.895000 1.615000 ;
        RECT 1.565000 1.075000 1.895000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.075000 1.345000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235000 0.275000 5.565000 0.725000 ;
        RECT 5.235000 0.725000 6.910000 0.905000 ;
        RECT 5.275000 1.785000 6.365000 1.955000 ;
        RECT 5.275000 1.955000 5.525000 2.465000 ;
        RECT 6.075000 0.275000 6.405000 0.725000 ;
        RECT 6.115000 1.415000 6.910000 1.655000 ;
        RECT 6.115000 1.655000 6.365000 1.785000 ;
        RECT 6.115000 1.955000 6.365000 2.465000 ;
        RECT 6.605000 0.905000 6.910000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.095000  0.255000 0.425000 0.725000 ;
      RECT 0.095000  0.725000 1.265000 0.735000 ;
      RECT 0.095000  0.735000 2.025000 0.905000 ;
      RECT 0.140000  1.795000 0.345000 2.635000 ;
      RECT 0.555000  1.785000 0.805000 2.295000 ;
      RECT 0.555000  2.295000 1.645000 2.465000 ;
      RECT 0.595000  0.085000 0.765000 0.555000 ;
      RECT 0.935000  0.255000 1.265000 0.725000 ;
      RECT 0.975000  1.785000 2.615000 1.955000 ;
      RECT 0.975000  1.955000 1.225000 2.125000 ;
      RECT 1.395000  2.125000 1.645000 2.295000 ;
      RECT 1.435000  0.085000 1.605000 0.555000 ;
      RECT 1.775000  0.255000 2.945000 0.475000 ;
      RECT 1.775000  0.475000 2.025000 0.735000 ;
      RECT 1.815000  2.125000 2.065000 2.635000 ;
      RECT 2.065000  1.075000 2.445000 1.415000 ;
      RECT 2.065000  1.415000 2.615000 1.785000 ;
      RECT 2.195000  0.645000 2.525000 0.815000 ;
      RECT 2.195000  0.815000 2.445000 1.075000 ;
      RECT 2.235000  1.955000 2.615000 1.965000 ;
      RECT 2.235000  1.965000 2.525000 2.465000 ;
      RECT 2.615000  1.075000 3.145000 1.245000 ;
      RECT 2.695000  2.135000 3.425000 2.635000 ;
      RECT 2.955000  0.725000 4.305000 0.905000 ;
      RECT 2.955000  0.905000 3.145000 1.075000 ;
      RECT 2.955000  1.245000 3.145000 1.785000 ;
      RECT 2.955000  1.785000 4.685000 1.965000 ;
      RECT 3.215000  0.085000 3.385000 0.555000 ;
      RECT 3.555000  0.305000 4.725000 0.475000 ;
      RECT 3.595000  1.965000 3.845000 2.125000 ;
      RECT 3.975000  0.645000 4.305000 0.725000 ;
      RECT 4.015000  2.135000 4.265000 2.635000 ;
      RECT 4.435000  1.965000 4.685000 2.465000 ;
      RECT 4.475000  0.475000 4.725000 0.895000 ;
      RECT 4.855000  1.795000 5.105000 2.635000 ;
      RECT 4.895000  0.085000 5.065000 0.895000 ;
      RECT 5.165000  1.075000 6.435000 1.245000 ;
      RECT 5.165000  1.245000 5.455000 1.615000 ;
      RECT 5.695000  2.165000 5.945000 2.635000 ;
      RECT 5.735000  0.085000 5.905000 0.555000 ;
      RECT 6.535000  1.825000 6.785000 2.635000 ;
      RECT 6.575000  0.085000 6.745000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.445000 2.615000 1.615000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.225000  1.445000 5.395000 1.615000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 2.385000 1.415000 2.675000 1.460000 ;
      RECT 2.385000 1.460000 5.455000 1.600000 ;
      RECT 2.385000 1.600000 2.675000 1.645000 ;
      RECT 5.165000 1.415000 5.455000 1.460000 ;
      RECT 5.165000 1.600000 5.455000 1.645000 ;
  END
END sky130_fd_sc_hd__o2bb2a_4
MACRO sky130_fd_sc_hd__o2bb2a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.770000 1.075000 1.220000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 0.380000 1.290000 0.735000 ;
        RECT 1.070000 0.735000 1.565000 0.905000 ;
        RECT 1.390000 0.905000 1.565000 1.100000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.250000 1.075000 3.595000 1.645000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.520000 1.075000 3.080000 1.325000 ;
        RECT 2.905000 1.325000 3.080000 2.425000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 0.825000 ;
        RECT 0.085000 0.825000 0.260000 1.795000 ;
        RECT 0.085000 1.795000 0.345000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.430000  0.995000 0.600000 1.445000 ;
      RECT 0.430000  1.445000 0.825000 1.615000 ;
      RECT 0.515000  2.235000 0.845000 2.635000 ;
      RECT 0.620000  0.085000 0.790000 0.750000 ;
      RECT 0.655000  1.615000 0.825000 1.885000 ;
      RECT 0.655000  1.885000 2.735000 2.055000 ;
      RECT 0.995000  1.495000 2.010000 1.715000 ;
      RECT 1.460000  0.395000 1.905000 0.565000 ;
      RECT 1.715000  2.235000 2.115000 2.635000 ;
      RECT 1.735000  0.565000 1.905000 1.355000 ;
      RECT 1.735000  1.355000 2.010000 1.495000 ;
      RECT 2.075000  0.320000 2.325000 0.690000 ;
      RECT 2.155000  0.690000 2.325000 1.075000 ;
      RECT 2.155000  1.075000 2.350000 1.245000 ;
      RECT 2.180000  1.245000 2.350000 1.495000 ;
      RECT 2.180000  1.495000 2.735000 1.885000 ;
      RECT 2.405000  2.055000 2.735000 2.290000 ;
      RECT 2.495000  0.320000 2.745000 0.725000 ;
      RECT 2.495000  0.725000 3.595000 0.905000 ;
      RECT 2.915000  0.085000 3.085000 0.555000 ;
      RECT 3.250000  1.815000 3.595000 2.635000 ;
      RECT 3.255000  0.320000 3.595000 0.725000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o2bb2a_1
MACRO sky130_fd_sc_hd__o2bb2a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.215000 1.075000 1.685000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 0.380000 1.735000 0.735000 ;
        RECT 1.515000 0.735000 2.020000 0.770000 ;
        RECT 1.515000 0.770000 2.025000 0.905000 ;
        RECT 1.855000 0.905000 2.025000 1.100000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.700000 1.075000 4.045000 1.645000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.075000 3.525000 1.325000 ;
        RECT 3.355000 1.325000 3.525000 2.425000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.870000 0.825000 ;
        RECT 0.535000 0.825000 0.705000 1.795000 ;
        RECT 0.535000 1.795000 0.790000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.135000 -0.085000 0.305000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.110000  0.085000 0.365000 0.910000 ;
      RECT 0.110000  1.410000 0.365000 2.635000 ;
      RECT 0.875000  0.995000 1.045000 1.445000 ;
      RECT 0.875000  1.445000 1.270000 1.615000 ;
      RECT 0.960000  2.235000 1.290000 2.635000 ;
      RECT 1.065000  0.085000 1.235000 0.750000 ;
      RECT 1.100000  1.615000 1.270000 1.885000 ;
      RECT 1.100000  1.885000 3.185000 2.055000 ;
      RECT 1.440000  1.495000 2.460000 1.715000 ;
      RECT 1.905000  0.395000 2.365000 0.565000 ;
      RECT 2.160000  2.235000 2.565000 2.635000 ;
      RECT 2.195000  0.565000 2.365000 1.355000 ;
      RECT 2.195000  1.355000 2.460000 1.495000 ;
      RECT 2.535000  0.320000 2.780000 0.690000 ;
      RECT 2.610000  0.690000 2.780000 1.075000 ;
      RECT 2.610000  1.075000 2.800000 1.245000 ;
      RECT 2.630000  1.245000 2.800000 1.495000 ;
      RECT 2.630000  1.495000 3.185000 1.885000 ;
      RECT 2.835000  2.055000 3.185000 2.425000 ;
      RECT 2.955000  0.320000 3.185000 0.725000 ;
      RECT 2.955000  0.725000 4.045000 0.905000 ;
      RECT 3.375000  0.085000 3.545000 0.555000 ;
      RECT 3.715000  0.320000 4.045000 0.725000 ;
      RECT 3.730000  1.815000 4.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o2bb2a_2
MACRO sky130_fd_sc_hd__dlygate4sd3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.775000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.210000 0.255000 3.595000 0.825000 ;
        RECT 3.210000 1.495000 3.595000 2.465000 ;
        RECT 3.315000 0.825000 3.595000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.200000  0.255000 0.485000 0.715000 ;
      RECT 0.200000  0.715000 1.155000 0.885000 ;
      RECT 0.200000  1.785000 1.155000 2.005000 ;
      RECT 0.200000  2.005000 0.485000 2.465000 ;
      RECT 0.655000  0.085000 0.925000 0.545000 ;
      RECT 0.655000  2.175000 0.925000 2.635000 ;
      RECT 0.945000  0.885000 1.155000 1.785000 ;
      RECT 1.325000  0.255000 1.725000 1.055000 ;
      RECT 1.325000  1.055000 2.420000 1.615000 ;
      RECT 1.325000  1.615000 1.725000 2.465000 ;
      RECT 1.915000  0.255000 2.195000 0.715000 ;
      RECT 1.915000  0.715000 3.040000 0.885000 ;
      RECT 1.915000  1.785000 3.040000 2.005000 ;
      RECT 1.915000  2.005000 2.195000 2.465000 ;
      RECT 2.590000  0.885000 3.040000 0.995000 ;
      RECT 2.590000  0.995000 3.145000 1.325000 ;
      RECT 2.590000  1.325000 3.040000 1.785000 ;
      RECT 2.715000  0.085000 3.040000 0.545000 ;
      RECT 2.715000  2.175000 3.040000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__dlygate4sd3_1
MACRO sky130_fd_sc_hd__a32oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775000 1.075000 5.465000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095000 1.075000 7.695000 1.300000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.295000 1.075000 9.985000 1.280000 ;
        RECT 9.805000 0.755000 9.985000 1.075000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.585000 0.995000 3.555000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.750000 1.305000 ;
        RECT 0.110000 1.305000 0.330000 1.965000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.575000 3.365000 1.745000 ;
        RECT 0.515000 1.745000 0.845000 2.085000 ;
        RECT 1.355000 1.745000 1.685000 2.085000 ;
        RECT 1.975000 0.990000 2.365000 1.575000 ;
        RECT 1.975000 1.745000 2.525000 2.085000 ;
        RECT 2.195000 0.635000 5.565000 0.805000 ;
        RECT 2.195000 0.805000 2.365000 0.990000 ;
        RECT 3.035000 1.745000 3.365000 2.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.095000  2.255000  3.705000 2.425000 ;
      RECT 0.175000  0.255000  0.345000 0.635000 ;
      RECT 0.175000  0.635000  2.025000 0.805000 ;
      RECT 0.515000  0.085000  0.845000 0.465000 ;
      RECT 1.015000  0.255000  1.185000 0.635000 ;
      RECT 1.355000  0.085000  1.685000 0.465000 ;
      RECT 1.855000  0.295000  3.785000 0.465000 ;
      RECT 1.855000  0.465000  2.025000 0.635000 ;
      RECT 3.535000  1.575000  9.925000 1.745000 ;
      RECT 3.535000  1.745000  3.705000 2.255000 ;
      RECT 3.895000  1.915000  4.225000 2.635000 ;
      RECT 3.975000  0.295000  7.805000 0.465000 ;
      RECT 4.395000  1.745000  4.565000 2.465000 ;
      RECT 4.770000  1.915000  5.440000 2.635000 ;
      RECT 5.640000  1.745000  5.810000 2.465000 ;
      RECT 6.215000  0.635000  9.505000 0.805000 ;
      RECT 6.215000  1.915000  6.545000 2.635000 ;
      RECT 6.715000  1.745000  6.885000 2.465000 ;
      RECT 7.055000  1.915000  7.385000 2.635000 ;
      RECT 7.555000  1.745000  7.725000 2.465000 ;
      RECT 7.995000  0.085000  8.325000 0.465000 ;
      RECT 8.415000  1.915000  8.745000 2.635000 ;
      RECT 8.495000  0.255000  8.665000 0.635000 ;
      RECT 8.835000  0.085000  9.165000 0.465000 ;
      RECT 8.915000  1.745000  9.085000 2.465000 ;
      RECT 9.255000  1.915000  9.585000 2.635000 ;
      RECT 9.335000  0.255000  9.505000 0.635000 ;
      RECT 9.685000  0.085000 10.025000 0.465000 ;
      RECT 9.755000  1.745000  9.925000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__a32oi_4
MACRO sky130_fd_sc_hd__a32oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.230000 1.075000 1.595000 1.255000 ;
        RECT 1.405000 0.345000 1.705000 0.765000 ;
        RECT 1.405000 0.765000 1.595000 1.075000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 0.995000 2.165000 1.325000 ;
        RECT 1.965000 0.415000 2.165000 0.995000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335000 1.015000 2.750000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 0.995000 1.025000 1.425000 ;
        RECT 0.855000 1.425000 1.255000 1.615000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.345000 1.325000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.575500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 1.165000 0.805000 ;
        RECT 0.515000 0.805000 0.685000 1.785000 ;
        RECT 0.515000 1.785000 0.865000 2.085000 ;
        RECT 0.915000 0.295000 1.165000 0.635000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.835000 0.345000 2.255000 ;
      RECT 0.085000  2.255000 1.345000 2.465000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 1.095000  1.785000 2.185000 1.955000 ;
      RECT 1.095000  1.955000 1.345000 2.255000 ;
      RECT 1.555000  2.135000 1.805000 2.635000 ;
      RECT 2.015000  1.745000 2.185000 1.785000 ;
      RECT 2.015000  1.955000 2.185000 2.465000 ;
      RECT 2.355000  0.085000 2.695000 0.805000 ;
      RECT 2.355000  1.495000 2.695000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a32oi_1
MACRO sky130_fd_sc_hd__a32oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415000 1.075000 3.220000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.075000 4.480000 1.625000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.715000 1.075000 5.860000 1.625000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.080000 1.725000 1.285000 ;
        RECT 1.175000 1.075000 1.505000 1.080000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.075000 0.825000 1.285000 ;
        RECT 0.145000 1.285000 0.325000 1.625000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.955000 0.845000 2.125000 ;
        RECT 0.595000 1.455000 2.180000 1.625000 ;
        RECT 0.595000 1.625000 0.765000 1.955000 ;
        RECT 1.355000 0.655000 3.100000 0.825000 ;
        RECT 1.435000 1.625000 1.605000 2.125000 ;
        RECT 1.965000 0.825000 2.180000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.095000  0.295000 0.425000 0.465000 ;
      RECT 0.175000  0.465000 0.345000 0.715000 ;
      RECT 0.175000  0.715000 1.185000 0.885000 ;
      RECT 0.175000  1.795000 0.345000 2.295000 ;
      RECT 0.175000  2.295000 2.025000 2.465000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 0.935000  0.295000 2.115000 0.465000 ;
      RECT 1.015000  0.465000 1.185000 0.715000 ;
      RECT 1.015000  1.795000 1.185000 2.295000 ;
      RECT 1.855000  1.795000 2.025000 1.915000 ;
      RECT 1.855000  1.915000 5.805000 2.085000 ;
      RECT 1.855000  2.085000 2.025000 2.295000 ;
      RECT 2.270000  2.255000 2.940000 2.635000 ;
      RECT 2.350000  0.295000 4.370000 0.465000 ;
      RECT 3.180000  1.795000 3.350000 1.915000 ;
      RECT 3.180000  2.085000 3.350000 2.465000 ;
      RECT 3.550000  2.255000 4.220000 2.635000 ;
      RECT 3.620000  0.635000 5.390000 0.805000 ;
      RECT 4.390000  1.795000 4.560000 1.915000 ;
      RECT 4.390000  2.085000 4.560000 2.465000 ;
      RECT 4.555000  0.085000 4.890000 0.465000 ;
      RECT 4.765000  2.255000 5.435000 2.635000 ;
      RECT 5.060000  0.275000 5.390000 0.635000 ;
      RECT 5.560000  0.085000 5.885000 0.885000 ;
      RECT 5.635000  1.795000 5.805000 1.915000 ;
      RECT 5.635000  2.085000 5.805000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__a32oi_2
MACRO sky130_fd_sc_hd__o311a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 0.995000 1.750000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.920000 0.995000 2.250000 1.325000 ;
        RECT 1.980000 1.325000 2.250000 2.070000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 0.995000 2.730000 1.325000 ;
        RECT 2.440000 1.325000 2.675000 2.070000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.900000 0.995000 3.300000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.810000 0.995000 4.055000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.905000 1.315000 ;
        RECT 0.550000 0.255000 0.825000 0.995000 ;
        RECT 0.550000 0.995000 0.905000 1.055000 ;
        RECT 0.550000 1.315000 0.905000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.085000 0.380000 0.885000 ;
      RECT 0.085000  1.485000 0.380000 2.635000 ;
      RECT 0.995000  0.085000 1.665000 0.825000 ;
      RECT 1.075000  0.995000 1.245000 1.495000 ;
      RECT 1.075000  1.495000 1.810000 1.665000 ;
      RECT 1.075000  1.835000 1.470000 2.635000 ;
      RECT 1.640000  1.665000 1.810000 2.295000 ;
      RECT 1.640000  2.295000 3.175000 2.465000 ;
      RECT 1.835000  0.310000 2.120000 0.655000 ;
      RECT 1.835000  0.655000 3.220000 0.825000 ;
      RECT 2.300000  0.085000 2.675000 0.485000 ;
      RECT 2.845000  1.495000 4.055000 1.665000 ;
      RECT 2.845000  1.665000 3.175000 2.295000 ;
      RECT 2.890000  0.310000 3.220000 0.655000 ;
      RECT 3.360000  1.835000 3.595000 2.635000 ;
      RECT 3.470000  0.255000 4.055000 0.825000 ;
      RECT 3.470000  0.825000 3.640000 1.495000 ;
      RECT 3.765000  1.665000 4.055000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o311a_2
MACRO sky130_fd_sc_hd__o311a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.995000 1.280000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.450000 0.995000 1.790000 1.325000 ;
        RECT 1.520000 1.325000 1.790000 2.070000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.980000 0.995000 2.270000 1.325000 ;
        RECT 1.980000 1.325000 2.215000 2.070000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 0.995000 2.840000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 0.995000 3.595000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.355000 1.070000 ;
        RECT 0.085000 1.070000 0.435000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.525000  0.085000 1.195000 0.825000 ;
      RECT 0.605000  0.995000 0.775000 1.495000 ;
      RECT 0.605000  1.495000 1.350000 1.665000 ;
      RECT 0.605000  1.835000 1.010000 2.635000 ;
      RECT 1.180000  1.665000 1.350000 2.295000 ;
      RECT 1.180000  2.295000 2.715000 2.465000 ;
      RECT 1.365000  0.310000 1.660000 0.655000 ;
      RECT 1.365000  0.655000 2.760000 0.825000 ;
      RECT 1.840000  0.085000 2.215000 0.485000 ;
      RECT 2.385000  1.495000 3.595000 1.665000 ;
      RECT 2.385000  1.665000 2.715000 2.295000 ;
      RECT 2.430000  0.310000 2.760000 0.655000 ;
      RECT 2.900000  1.835000 3.135000 2.635000 ;
      RECT 3.010000  0.255000 3.595000 0.825000 ;
      RECT 3.010000  0.825000 3.180000 1.495000 ;
      RECT 3.305000  1.665000 3.595000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o311a_1
MACRO sky130_fd_sc_hd__o311a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.950000 1.055000 7.735000 1.315000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.020000 1.055000 6.770000 1.315000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.655000 1.055000 5.850000 1.315000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.250000 1.055000 4.475000 1.315000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.115000 1.055000 3.080000 1.315000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.765000 1.315000 ;
        RECT 0.595000 0.255000 0.765000 0.715000 ;
        RECT 0.595000 0.715000 1.605000 0.885000 ;
        RECT 0.595000 0.885000 0.765000 1.055000 ;
        RECT 0.595000 1.315000 0.765000 1.485000 ;
        RECT 0.595000 1.485000 1.605000 1.725000 ;
        RECT 0.595000 1.725000 0.765000 2.465000 ;
        RECT 1.435000 0.255000 1.605000 0.715000 ;
        RECT 1.435000 1.725000 1.605000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.085000 0.425000 0.885000 ;
      RECT 0.085000  1.485000 0.425000 2.635000 ;
      RECT 0.935000  0.085000 1.265000 0.545000 ;
      RECT 0.935000  1.055000 1.945000 1.315000 ;
      RECT 0.935000  1.895000 1.265000 2.635000 ;
      RECT 1.775000  0.085000 2.025000 0.545000 ;
      RECT 1.775000  0.715000 3.045000 0.885000 ;
      RECT 1.775000  0.885000 1.945000 1.055000 ;
      RECT 1.775000  1.315000 1.945000 1.485000 ;
      RECT 1.775000  1.485000 5.005000 1.725000 ;
      RECT 1.775000  1.895000 2.445000 2.635000 ;
      RECT 2.195000  0.255000 4.305000 0.505000 ;
      RECT 2.195000  0.675000 3.045000 0.715000 ;
      RECT 2.615000  1.725000 2.785000 2.465000 ;
      RECT 2.955000  1.895000 3.285000 2.635000 ;
      RECT 3.215000  0.505000 3.385000 0.885000 ;
      RECT 3.455000  1.725000 3.625000 2.465000 ;
      RECT 3.555000  0.675000 7.735000 0.885000 ;
      RECT 3.855000  1.895000 4.045000 2.635000 ;
      RECT 4.335000  1.895000 4.665000 2.295000 ;
      RECT 4.335000  2.295000 6.445000 2.465000 ;
      RECT 4.485000  0.255000 4.755000 0.675000 ;
      RECT 4.835000  1.725000 5.005000 2.125000 ;
      RECT 4.925000  0.085000 5.605000 0.505000 ;
      RECT 5.255000  1.485000 5.525000 2.295000 ;
      RECT 5.695000  1.485000 7.735000 1.725000 ;
      RECT 5.695000  1.725000 5.945000 2.125000 ;
      RECT 5.775000  0.255000 5.945000 0.675000 ;
      RECT 6.115000  0.085000 6.445000 0.505000 ;
      RECT 6.115000  1.895000 6.445000 2.295000 ;
      RECT 6.615000  0.255000 6.785000 0.675000 ;
      RECT 6.615000  1.725000 6.785000 2.125000 ;
      RECT 6.955000  0.085000 7.285000 0.505000 ;
      RECT 6.955000  1.895000 7.285000 2.635000 ;
      RECT 7.455000  0.255000 7.735000 0.675000 ;
      RECT 7.455000  1.725000 7.735000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__o311a_4
MACRO sky130_fd_sc_hd__o21bai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21bai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195000 1.075000 2.675000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.075000 2.025000 1.285000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.535000 1.345000 ;
        RECT 0.085000 1.345000 0.355000 2.445000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.474000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 0.255000 1.285000 0.645000 ;
        RECT 1.115000 0.645000 1.355000 0.825000 ;
        RECT 1.185000 0.825000 1.355000 1.455000 ;
        RECT 1.185000 1.455000 1.795000 1.625000 ;
        RECT 1.470000 1.625000 1.795000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.085000 0.360000 0.825000 ;
      RECT 0.525000  1.535000 1.015000 1.705000 ;
      RECT 0.525000  1.705000 0.800000 2.210000 ;
      RECT 0.580000  0.495000 0.770000 0.655000 ;
      RECT 0.580000  0.655000 0.890000 0.825000 ;
      RECT 0.720000  0.825000 0.890000 0.995000 ;
      RECT 0.720000  0.995000 1.015000 1.535000 ;
      RECT 0.970000  1.875000 1.300000 2.635000 ;
      RECT 1.490000  0.255000 1.820000 0.485000 ;
      RECT 1.570000  0.485000 1.740000 0.735000 ;
      RECT 1.570000  0.735000 2.665000 0.905000 ;
      RECT 1.995000  0.085000 2.165000 0.555000 ;
      RECT 2.270000  1.535000 2.645000 2.635000 ;
      RECT 2.335000  0.270000 2.665000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__o21bai_1
MACRO sky130_fd_sc_hd__o21bai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21bai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.260000 1.075000 4.055000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.950000 1.075000 3.090000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.525000 1.325000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.445000 2.650000 1.615000 ;
        RECT 1.085000 1.615000 1.255000 2.465000 ;
        RECT 1.525000 0.645000 1.855000 0.905000 ;
        RECT 1.525000 0.905000 1.780000 1.445000 ;
        RECT 2.405000 1.615000 2.650000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.180000  0.085000 0.350000 0.825000 ;
      RECT 0.180000  1.495000 0.865000 1.665000 ;
      RECT 0.180000  1.665000 0.350000 1.915000 ;
      RECT 0.585000  1.875000 0.915000 2.635000 ;
      RECT 0.600000  0.445000 0.865000 0.825000 ;
      RECT 0.695000  0.825000 0.865000 1.075000 ;
      RECT 0.695000  1.075000 1.335000 1.245000 ;
      RECT 0.695000  1.245000 0.865000 1.495000 ;
      RECT 1.075000  0.255000 2.275000 0.475000 ;
      RECT 1.075000  0.475000 1.355000 0.905000 ;
      RECT 1.470000  1.795000 1.720000 2.635000 ;
      RECT 1.955000  1.795000 2.235000 2.295000 ;
      RECT 1.955000  2.295000 3.035000 2.465000 ;
      RECT 2.025000  0.475000 2.275000 0.725000 ;
      RECT 2.025000  0.725000 3.980000 0.905000 ;
      RECT 2.445000  0.085000 2.615000 0.555000 ;
      RECT 2.785000  0.255000 3.115000 0.725000 ;
      RECT 2.865000  1.455000 3.980000 1.665000 ;
      RECT 2.865000  1.665000 3.035000 2.295000 ;
      RECT 3.205000  1.835000 3.535000 2.635000 ;
      RECT 3.285000  0.085000 3.455000 0.555000 ;
      RECT 3.625000  0.265000 3.980000 0.725000 ;
      RECT 3.705000  1.665000 3.980000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o21bai_2
MACRO sky130_fd_sc_hd__o21bai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21bai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.645000 1.075000 6.810000 1.285000 ;
        RECT 6.585000 1.285000 6.810000 2.455000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.065000 1.075000 4.475000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.555000 1.285000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.455000 4.315000 1.625000 ;
        RECT 1.065000 1.625000 1.275000 2.465000 ;
        RECT 1.420000 0.645000 2.675000 0.815000 ;
        RECT 1.865000 1.625000 2.115000 2.465000 ;
        RECT 2.445000 0.815000 2.675000 1.075000 ;
        RECT 2.445000 1.075000 2.895000 1.445000 ;
        RECT 2.445000 1.445000 4.315000 1.455000 ;
        RECT 3.225000 1.625000 3.475000 2.125000 ;
        RECT 4.065000 1.625000 4.315000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.145000  1.455000 0.895000 1.625000 ;
      RECT 0.145000  1.625000 0.475000 2.435000 ;
      RECT 0.225000  0.085000 0.395000 0.895000 ;
      RECT 0.565000  0.290000 0.895000 0.895000 ;
      RECT 0.645000  1.795000 0.855000 2.635000 ;
      RECT 0.725000  0.895000 0.895000 1.075000 ;
      RECT 0.725000  1.075000 2.275000 1.285000 ;
      RECT 0.725000  1.285000 0.895000 1.455000 ;
      RECT 1.080000  0.305000 3.095000 0.475000 ;
      RECT 1.445000  1.795000 1.695000 2.635000 ;
      RECT 2.285000  1.795000 2.535000 2.635000 ;
      RECT 2.775000  1.795000 3.055000 2.295000 ;
      RECT 2.775000  2.295000 4.735000 2.465000 ;
      RECT 2.845000  0.475000 3.095000 0.725000 ;
      RECT 2.845000  0.725000 6.455000 0.905000 ;
      RECT 3.265000  0.085000 3.435000 0.555000 ;
      RECT 3.605000  0.255000 3.935000 0.725000 ;
      RECT 3.645000  1.795000 3.895000 2.295000 ;
      RECT 4.105000  0.085000 4.275000 0.555000 ;
      RECT 4.445000  0.255000 4.775000 0.725000 ;
      RECT 4.485000  1.455000 6.415000 1.625000 ;
      RECT 4.485000  1.625000 4.735000 2.295000 ;
      RECT 4.905000  1.795000 5.155000 2.635000 ;
      RECT 4.945000  0.085000 5.115000 0.555000 ;
      RECT 5.285000  0.255000 5.615000 0.725000 ;
      RECT 5.325000  1.625000 5.575000 2.465000 ;
      RECT 5.745000  1.795000 5.995000 2.635000 ;
      RECT 5.785000  0.085000 5.955000 0.555000 ;
      RECT 6.125000  0.255000 6.455000 0.725000 ;
      RECT 6.165000  1.625000 6.415000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
END sky130_fd_sc_hd__o21bai_4
MACRO sky130_fd_sc_hd__nor4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.115000 0.995000 3.595000 1.275000 ;
        RECT 3.295000 1.275000 3.595000 1.705000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615000 0.995000 2.945000 1.445000 ;
        RECT 2.615000 1.445000 3.085000 1.630000 ;
        RECT 2.825000 1.630000 3.085000 2.410000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.780000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.995000 1.240000 1.325000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.606900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.470000 1.955000 2.055000 2.125000 ;
        RECT 1.855000 0.655000 3.085000 0.825000 ;
        RECT 1.855000 0.825000 2.055000 1.955000 ;
        RECT 2.015000 0.300000 2.215000 0.655000 ;
        RECT 2.885000 0.310000 3.085000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.450000 0.405000 0.825000 ;
      RECT 0.085000  0.825000 0.260000 1.885000 ;
      RECT 0.085000  1.885000 1.205000 2.070000 ;
      RECT 0.085000  2.070000 0.345000 2.455000 ;
      RECT 0.515000  2.240000 0.845000 2.635000 ;
      RECT 0.655000  0.085000 0.825000 0.825000 ;
      RECT 0.995000  1.525000 1.590000 1.715000 ;
      RECT 1.035000  2.070000 1.205000 2.295000 ;
      RECT 1.035000  2.295000 2.395000 2.465000 ;
      RECT 1.075000  0.450000 1.245000 0.655000 ;
      RECT 1.075000  0.655000 1.590000 0.825000 ;
      RECT 1.410000  0.825000 1.590000 0.995000 ;
      RECT 1.410000  0.995000 1.685000 1.325000 ;
      RECT 1.410000  1.325000 1.590000 1.525000 ;
      RECT 1.515000  0.085000 1.845000 0.480000 ;
      RECT 2.225000  0.995000 2.395000 2.295000 ;
      RECT 2.385000  0.085000 2.715000 0.485000 ;
      RECT 3.255000  0.085000 3.585000 0.825000 ;
      RECT 3.255000  1.875000 3.585000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4bb_1
MACRO sky130_fd_sc_hd__nor4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.375000 1.075000 9.110000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.150000 1.075000 7.105000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.445000 1.365000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.075000 1.295000 1.325000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.840000 1.415000 3.185000 1.705000 ;
        RECT 1.935000 0.255000 2.265000 0.725000 ;
        RECT 1.935000 0.725000 8.665000 0.905000 ;
        RECT 2.775000 0.255000 3.105000 0.725000 ;
        RECT 3.015000 0.905000 3.185000 1.415000 ;
        RECT 3.615000 0.255000 3.945000 0.725000 ;
        RECT 4.455000 0.255000 4.785000 0.725000 ;
        RECT 5.815000 0.255000 6.145000 0.725000 ;
        RECT 6.655000 0.255000 6.985000 0.725000 ;
        RECT 7.495000 0.255000 7.825000 0.725000 ;
        RECT 8.335000 0.255000 8.665000 0.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.085000  0.255000 0.445000 0.725000 ;
      RECT 0.085000  0.725000 0.785000 0.895000 ;
      RECT 0.085000  1.535000 0.785000 1.875000 ;
      RECT 0.085000  1.875000 3.525000 2.045000 ;
      RECT 0.085000  2.045000 0.365000 2.465000 ;
      RECT 0.535000  2.215000 0.865000 2.635000 ;
      RECT 0.615000  0.085000 0.785000 0.555000 ;
      RECT 0.615000  0.895000 0.785000 1.535000 ;
      RECT 0.955000  0.255000 1.285000 0.735000 ;
      RECT 0.955000  0.735000 1.635000 0.905000 ;
      RECT 0.955000  1.535000 1.635000 1.705000 ;
      RECT 1.465000  0.905000 1.635000 1.075000 ;
      RECT 1.465000  1.075000 2.845000 1.245000 ;
      RECT 1.465000  1.245000 1.635000 1.535000 ;
      RECT 1.515000  2.215000 3.525000 2.295000 ;
      RECT 1.515000  2.295000 5.195000 2.465000 ;
      RECT 1.595000  0.085000 1.765000 0.555000 ;
      RECT 2.435000  0.085000 2.605000 0.555000 ;
      RECT 3.275000  0.085000 3.445000 0.555000 ;
      RECT 3.355000  1.075000 4.905000 1.285000 ;
      RECT 3.355000  1.285000 3.525000 1.875000 ;
      RECT 3.695000  1.455000 6.945000 1.625000 ;
      RECT 3.695000  1.625000 3.905000 2.125000 ;
      RECT 4.075000  1.795000 4.325000 2.295000 ;
      RECT 4.115000  0.085000 4.285000 0.555000 ;
      RECT 4.495000  1.625000 4.745000 2.125000 ;
      RECT 4.915000  1.795000 5.195000 2.295000 ;
      RECT 4.955000  0.085000 5.645000 0.555000 ;
      RECT 5.380000  1.795000 5.685000 2.295000 ;
      RECT 5.380000  2.295000 7.365000 2.465000 ;
      RECT 5.855000  1.625000 6.105000 2.125000 ;
      RECT 6.275000  1.795000 6.525000 2.295000 ;
      RECT 6.315000  0.085000 6.485000 0.555000 ;
      RECT 6.695000  1.625000 6.945000 2.125000 ;
      RECT 7.115000  1.455000 9.110000 1.625000 ;
      RECT 7.115000  1.625000 7.365000 2.295000 ;
      RECT 7.155000  0.085000 7.325000 0.555000 ;
      RECT 7.535000  1.795000 7.785000 2.635000 ;
      RECT 7.955000  1.625000 8.205000 2.465000 ;
      RECT 7.995000  0.085000 8.165000 0.555000 ;
      RECT 8.375000  1.795000 8.625000 2.635000 ;
      RECT 8.795000  1.625000 9.110000 2.465000 ;
      RECT 8.835000  0.085000 9.110000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4bb_4
MACRO sky130_fd_sc_hd__nor4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.130000 1.075000 5.895000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 1.075000 4.960000 1.275000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.995000 1.235000 1.325000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.780000 1.695000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.060000 0.255000 2.390000 0.725000 ;
        RECT 2.060000 0.725000 5.450000 0.905000 ;
        RECT 2.900000 0.255000 3.230000 0.725000 ;
        RECT 2.900000 1.445000 3.995000 1.705000 ;
        RECT 3.575000 0.905000 3.995000 1.445000 ;
        RECT 4.280000 0.255000 4.610000 0.725000 ;
        RECT 5.120000 0.255000 5.450000 0.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.450000 0.465000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.885000 ;
      RECT 0.085000  1.885000 1.915000 2.055000 ;
      RECT 0.085000  2.055000 0.345000 2.455000 ;
      RECT 0.515000  2.240000 0.845000 2.635000 ;
      RECT 0.635000  0.085000 0.805000 0.825000 ;
      RECT 0.995000  1.525000 1.575000 1.715000 ;
      RECT 1.055000  0.450000 1.250000 0.655000 ;
      RECT 1.055000  0.655000 1.575000 0.825000 ;
      RECT 1.405000  0.825000 1.575000 1.075000 ;
      RECT 1.405000  1.075000 2.390000 1.245000 ;
      RECT 1.405000  1.245000 1.575000 1.525000 ;
      RECT 1.560000  0.085000 1.890000 0.480000 ;
      RECT 1.640000  2.225000 1.970000 2.295000 ;
      RECT 1.640000  2.295000 3.650000 2.465000 ;
      RECT 1.745000  1.415000 2.730000 1.585000 ;
      RECT 1.745000  1.585000 1.915000 1.885000 ;
      RECT 2.140000  1.795000 2.310000 1.875000 ;
      RECT 2.140000  1.875000 4.610000 2.045000 ;
      RECT 2.140000  2.045000 2.310000 2.125000 ;
      RECT 2.480000  2.215000 3.650000 2.295000 ;
      RECT 2.560000  0.085000 2.730000 0.555000 ;
      RECT 2.560000  1.075000 3.405000 1.275000 ;
      RECT 2.560000  1.275000 2.730000 1.415000 ;
      RECT 3.400000  0.085000 4.110000 0.555000 ;
      RECT 3.860000  2.215000 4.990000 2.465000 ;
      RECT 4.320000  1.455000 4.610000 1.875000 ;
      RECT 4.780000  0.085000 4.950000 0.555000 ;
      RECT 4.780000  1.455000 5.870000 1.625000 ;
      RECT 4.780000  1.625000 4.990000 2.215000 ;
      RECT 5.160000  1.795000 5.370000 2.635000 ;
      RECT 5.540000  1.625000 5.870000 2.465000 ;
      RECT 5.620000  0.085000 5.895000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4bb_2
MACRO sky130_fd_sc_hd__sdfbbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfbbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.26000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 1.325000 4.025000 2.375000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.915000 0.255000 14.175000 0.825000 ;
        RECT 13.915000 1.605000 14.175000 2.465000 ;
        RECT 13.965000 0.825000 14.175000 1.605000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.500000 0.255000 12.785000 0.715000 ;
        RECT 12.500000 1.630000 12.785000 2.465000 ;
        RECT 12.605000 0.715000 12.785000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.535000 1.095000 11.990000 1.325000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 1.025000 1.720000 1.685000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 0.345000 2.180000 0.845000 ;
        RECT 1.960000 0.845000 2.415000 1.015000 ;
        RECT 1.960000 1.015000 2.180000 1.695000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 0.735000 6.295000 0.965000 ;
        RECT 5.885000 0.965000 6.215000 1.065000 ;
      LAYER mcon ;
        RECT 6.125000 0.765000 6.295000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755000 0.735000 10.130000 1.065000 ;
      LAYER mcon ;
        RECT 9.805000 0.765000 9.975000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065000 0.735000  6.355000 0.780000 ;
        RECT 6.065000 0.780000 10.035000 0.920000 ;
        RECT 6.065000 0.920000  6.355000 0.965000 ;
        RECT 9.745000 0.735000 10.035000 0.780000 ;
        RECT 9.745000 0.920000 10.035000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 14.450000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.170000  0.345000  0.345000 0.635000 ;
      RECT  0.170000  0.635000  0.835000 0.805000 ;
      RECT  0.170000  1.795000  0.835000 1.965000 ;
      RECT  0.170000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.605000  0.805000  0.835000 1.795000 ;
      RECT  1.015000  0.345000  1.240000 2.465000 ;
      RECT  1.455000  0.085000  1.705000 0.635000 ;
      RECT  1.455000  1.885000  1.785000 2.635000 ;
      RECT  2.235000  1.875000  2.565000 2.385000 ;
      RECT  2.350000  0.265000  2.755000 0.595000 ;
      RECT  2.350000  1.185000  3.075000 1.365000 ;
      RECT  2.350000  1.365000  2.565000 1.875000 ;
      RECT  2.585000  0.595000  2.755000 1.075000 ;
      RECT  2.585000  1.075000  3.075000 1.185000 ;
      RECT  2.745000  1.575000  3.645000 1.745000 ;
      RECT  2.745000  1.745000  3.065000 1.905000 ;
      RECT  2.895000  1.905000  3.065000 2.465000 ;
      RECT  2.925000  0.305000  3.125000 0.625000 ;
      RECT  2.925000  0.625000  3.645000 0.765000 ;
      RECT  2.925000  0.765000  3.770000 0.795000 ;
      RECT  3.310000  2.215000  3.640000 2.635000 ;
      RECT  3.370000  0.085000  3.700000 0.445000 ;
      RECT  3.475000  0.795000  3.770000 1.095000 ;
      RECT  3.475000  1.095000  3.645000 1.575000 ;
      RECT  4.230000  0.305000  4.455000 2.465000 ;
      RECT  4.625000  0.705000  4.845000 1.575000 ;
      RECT  4.625000  1.575000  5.125000 1.955000 ;
      RECT  4.635000  2.250000  5.465000 2.420000 ;
      RECT  4.700000  0.265000  5.715000 0.465000 ;
      RECT  5.025000  0.645000  5.375000 1.015000 ;
      RECT  5.295000  1.195000  5.715000 1.235000 ;
      RECT  5.295000  1.235000  6.645000 1.405000 ;
      RECT  5.295000  1.405000  5.465000 2.250000 ;
      RECT  5.545000  0.465000  5.715000 1.195000 ;
      RECT  5.635000  1.575000  5.885000 1.785000 ;
      RECT  5.635000  1.785000  6.985000 2.035000 ;
      RECT  5.705000  2.205000  6.085000 2.635000 ;
      RECT  5.885000  0.085000  6.055000 0.525000 ;
      RECT  6.225000  0.255000  7.395000 0.425000 ;
      RECT  6.225000  0.425000  6.555000 0.465000 ;
      RECT  6.385000  2.035000  6.555000 2.375000 ;
      RECT  6.395000  1.405000  6.645000 1.485000 ;
      RECT  6.425000  1.155000  6.645000 1.235000 ;
      RECT  6.700000  0.595000  7.030000 0.765000 ;
      RECT  6.815000  0.765000  7.030000 0.895000 ;
      RECT  6.815000  0.895000  8.125000 1.065000 ;
      RECT  6.815000  1.065000  6.985000 1.785000 ;
      RECT  7.155000  1.235000  7.485000 1.415000 ;
      RECT  7.155000  1.415000  8.160000 1.655000 ;
      RECT  7.175000  1.915000  7.505000 2.635000 ;
      RECT  7.200000  0.425000  7.395000 0.715000 ;
      RECT  7.640000  0.085000  7.975000 0.465000 ;
      RECT  7.795000  1.065000  8.125000 1.235000 ;
      RECT  8.360000  1.575000  8.595000 1.985000 ;
      RECT  8.420000  0.705000  8.705000 1.125000 ;
      RECT  8.420000  1.125000  9.040000 1.305000 ;
      RECT  8.550000  2.250000  9.380000 2.420000 ;
      RECT  8.615000  0.265000  9.380000 0.465000 ;
      RECT  8.835000  1.305000  9.040000 1.905000 ;
      RECT  9.210000  0.465000  9.380000 1.235000 ;
      RECT  9.210000  1.235000 10.560000 1.405000 ;
      RECT  9.210000  1.405000  9.380000 2.250000 ;
      RECT  9.550000  1.575000  9.800000 1.915000 ;
      RECT  9.550000  1.915000 12.330000 2.085000 ;
      RECT  9.560000  0.085000  9.820000 0.525000 ;
      RECT  9.620000  2.255000 10.000000 2.635000 ;
      RECT 10.080000  0.255000 11.250000 0.425000 ;
      RECT 10.080000  0.425000 10.430000 0.465000 ;
      RECT 10.240000  2.085000 10.410000 2.375000 ;
      RECT 10.340000  1.075000 10.560000 1.235000 ;
      RECT 10.575000  0.645000 10.905000 0.815000 ;
      RECT 10.730000  0.815000 10.905000 1.915000 ;
      RECT 10.940000  2.255000 12.330000 2.635000 ;
      RECT 11.075000  0.425000 11.250000 0.585000 ;
      RECT 11.080000  0.755000 11.765000 0.925000 ;
      RECT 11.080000  0.925000 11.355000 1.575000 ;
      RECT 11.080000  1.575000 11.855000 1.745000 ;
      RECT 11.565000  0.265000 11.765000 0.755000 ;
      RECT 12.000000  0.085000 12.330000 0.805000 ;
      RECT 12.160000  0.995000 12.425000 1.325000 ;
      RECT 12.160000  1.325000 12.330000 1.915000 ;
      RECT 12.960000  0.255000 13.275000 0.995000 ;
      RECT 12.960000  0.995000 13.795000 1.325000 ;
      RECT 12.960000  1.325000 13.275000 2.415000 ;
      RECT 13.450000  1.765000 13.745000 2.635000 ;
      RECT 13.455000  0.085000 13.745000 0.545000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  1.785000  0.775000 1.955000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  0.765000  1.235000 0.935000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  1.105000  3.075000 1.275000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.785000  4.915000 1.955000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  0.765000  5.375000 0.935000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  1.445000  8.135000 1.615000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  1.105000  8.595000 1.275000 ;
      RECT  8.425000  1.785000  8.595000 1.955000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  1.445000 11.355000 1.615000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT  0.545000 1.755000  0.835000 1.800000 ;
      RECT  0.545000 1.800000  8.655000 1.940000 ;
      RECT  0.545000 1.940000  0.835000 1.985000 ;
      RECT  1.005000 0.735000  1.295000 0.780000 ;
      RECT  1.005000 0.780000  5.435000 0.920000 ;
      RECT  1.005000 0.920000  1.295000 0.965000 ;
      RECT  2.845000 1.075000  3.135000 1.120000 ;
      RECT  2.845000 1.120000  4.515000 1.260000 ;
      RECT  2.845000 1.260000  3.135000 1.305000 ;
      RECT  4.225000 1.075000  4.515000 1.120000 ;
      RECT  4.225000 1.260000  4.515000 1.305000 ;
      RECT  4.685000 1.755000  4.975000 1.800000 ;
      RECT  4.685000 1.940000  4.975000 1.985000 ;
      RECT  5.145000 0.735000  5.435000 0.780000 ;
      RECT  5.145000 0.920000  5.435000 0.965000 ;
      RECT  5.220000 0.965000  5.435000 1.120000 ;
      RECT  5.220000 1.120000  8.655000 1.260000 ;
      RECT  7.905000 1.415000  8.195000 1.460000 ;
      RECT  7.905000 1.460000 11.415000 1.600000 ;
      RECT  7.905000 1.600000  8.195000 1.645000 ;
      RECT  8.365000 1.075000  8.655000 1.120000 ;
      RECT  8.365000 1.260000  8.655000 1.305000 ;
      RECT  8.365000 1.755000  8.655000 1.800000 ;
      RECT  8.365000 1.940000  8.655000 1.985000 ;
      RECT 11.125000 1.415000 11.415000 1.460000 ;
      RECT 11.125000 1.600000 11.415000 1.645000 ;
  END
END sky130_fd_sc_hd__sdfbbp_1
MACRO sky130_fd_sc_hd__lpflow_inputiso0p_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso0p_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 1.645000 2.175000 1.955000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.445000 1.615000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.350000 1.580000 2.655000 2.365000 ;
        RECT 2.415000 0.255000 2.655000 0.775000 ;
        RECT 2.480000 0.775000 2.655000 1.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.590000 ;
      RECT 0.175000  1.785000 0.850000 2.015000 ;
      RECT 0.175000  2.015000 0.345000 2.445000 ;
      RECT 0.515000  2.185000 0.845000 2.635000 ;
      RECT 0.595000  0.280000 0.835000 0.655000 ;
      RECT 0.615000  0.655000 0.835000 0.805000 ;
      RECT 0.615000  0.805000 1.150000 1.135000 ;
      RECT 0.615000  1.135000 0.850000 1.785000 ;
      RECT 1.020000  1.305000 2.305000 1.325000 ;
      RECT 1.020000  1.325000 1.880000 1.475000 ;
      RECT 1.020000  1.475000 1.305000 2.420000 ;
      RECT 1.115000  0.270000 1.285000 0.415000 ;
      RECT 1.115000  0.415000 1.490000 0.610000 ;
      RECT 1.320000  0.610000 1.490000 0.945000 ;
      RECT 1.320000  0.945000 2.305000 1.305000 ;
      RECT 1.485000  2.165000 2.170000 2.635000 ;
      RECT 1.850000  0.085000 2.245000 0.580000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso0p_1
MACRO sky130_fd_sc_hd__o32ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.750000 1.075000 5.865000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.370000 1.075000 4.480000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.075000 3.065000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 1.075000 1.705000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.845000 1.325000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.655000 2.045000 0.905000 ;
        RECT 0.515000 1.495000 3.105000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.095000 ;
        RECT 1.875000 0.905000 2.045000 1.105000 ;
        RECT 1.875000 1.105000 2.170000 1.495000 ;
        RECT 2.775000 1.665000 3.105000 2.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.090000  0.255000 2.405000 0.485000 ;
      RECT 0.090000  0.485000 0.345000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.295000 ;
      RECT 0.090000  2.295000 1.265000 2.465000 ;
      RECT 1.015000  1.835000 2.105000 2.005000 ;
      RECT 1.015000  2.005000 1.265000 2.295000 ;
      RECT 1.435000  2.175000 1.605000 2.635000 ;
      RECT 1.775000  2.005000 2.105000 2.455000 ;
      RECT 2.235000  0.485000 2.405000 0.715000 ;
      RECT 2.235000  0.715000 5.755000 0.905000 ;
      RECT 2.335000  1.835000 2.585000 2.255000 ;
      RECT 2.335000  2.255000 4.385000 2.445000 ;
      RECT 2.620000  0.085000 2.950000 0.545000 ;
      RECT 3.135000  0.255000 3.465000 0.715000 ;
      RECT 3.275000  1.495000 3.445000 2.255000 ;
      RECT 3.615000  1.495000 5.325000 1.665000 ;
      RECT 3.615000  1.665000 3.945000 2.085000 ;
      RECT 3.635000  0.085000 3.805000 0.545000 ;
      RECT 4.055000  0.255000 4.725000 0.715000 ;
      RECT 4.135000  1.835000 4.385000 2.255000 ;
      RECT 4.620000  1.835000 4.825000 2.635000 ;
      RECT 4.905000  0.085000 5.235000 0.545000 ;
      RECT 4.995000  1.665000 5.325000 2.460000 ;
      RECT 5.425000  0.255000 5.755000 0.715000 ;
      RECT 5.495000  1.495000 5.715000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__o32ai_2
MACRO sky130_fd_sc_hd__o32ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.575000 0.995000 3.135000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.930000 0.995000 2.225000 2.465000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.410000 0.995000 1.700000 1.615000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.685000 0.345000 0.995000 ;
        RECT 0.090000 0.995000 0.360000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.870000 0.995000 1.240000 1.615000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.821250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.655000 0.845000 0.825000 ;
        RECT 0.530000 0.825000 0.700000 1.785000 ;
        RECT 0.530000 1.785000 1.545000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  0.255000 1.345000 0.485000 ;
      RECT 0.090000  1.495000 0.360000 2.635000 ;
      RECT 1.015000  0.485000 1.345000 0.655000 ;
      RECT 1.015000  0.655000 2.525000 0.825000 ;
      RECT 1.515000  0.085000 2.185000 0.485000 ;
      RECT 2.355000  0.375000 2.525000 0.655000 ;
      RECT 2.695000  0.085000 3.135000 0.825000 ;
      RECT 2.695000  1.495000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o32ai_1
MACRO sky130_fd_sc_hd__o32ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.290000 1.075000 10.035000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.090000 1.075000 7.260000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.770000 1.075000 5.380000 1.275000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.205000 1.075000 3.540000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.685000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.655000 3.380000 0.905000 ;
        RECT 0.515000 1.495000 5.580000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.085000 ;
        RECT 1.355000 1.665000 1.700000 2.085000 ;
        RECT 1.855000 0.905000 2.035000 1.495000 ;
        RECT 4.410000 1.665000 4.740000 2.085000 ;
        RECT 5.250000 1.665000 5.580000 2.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.090000  0.255000  3.800000 0.465000 ;
      RECT 0.090000  0.465000  0.345000 0.905000 ;
      RECT 0.090000  1.495000  0.345000 2.255000 ;
      RECT 0.090000  2.255000  2.040000 2.465000 ;
      RECT 1.015000  1.835000  1.185000 2.255000 ;
      RECT 1.870000  1.835000  3.800000 2.005000 ;
      RECT 1.870000  2.005000  2.040000 2.255000 ;
      RECT 2.210000  2.175000  2.540000 2.635000 ;
      RECT 2.710000  2.005000  2.880000 2.425000 ;
      RECT 3.050000  2.175000  3.380000 2.635000 ;
      RECT 3.550000  0.465000  3.800000 0.735000 ;
      RECT 3.550000  0.735000 10.035000 0.905000 ;
      RECT 3.550000  2.005000  3.800000 2.465000 ;
      RECT 3.970000  0.085000  4.140000 0.545000 ;
      RECT 3.990000  1.835000  4.240000 2.255000 ;
      RECT 3.990000  2.255000  7.680000 2.465000 ;
      RECT 4.310000  0.255000  4.640000 0.735000 ;
      RECT 4.810000  0.085000  5.140000 0.545000 ;
      RECT 4.910000  1.835000  5.080000 2.255000 ;
      RECT 5.310000  0.255000  5.980000 0.735000 ;
      RECT 5.750000  1.835000  5.920000 2.255000 ;
      RECT 6.090000  1.495000  9.460000 1.665000 ;
      RECT 6.090000  1.665000  6.420000 2.085000 ;
      RECT 6.170000  0.085000  6.340000 0.545000 ;
      RECT 6.510000  0.255000  6.840000 0.735000 ;
      RECT 6.590000  1.835000  6.760000 2.255000 ;
      RECT 6.930000  1.665000  7.260000 2.085000 ;
      RECT 7.010000  0.085000  7.180000 0.545000 ;
      RECT 7.350000  0.255000  8.040000 0.735000 ;
      RECT 7.430000  1.835000  7.680000 2.255000 ;
      RECT 7.870000  1.835000  8.120000 2.635000 ;
      RECT 8.290000  1.665000  8.620000 2.465000 ;
      RECT 8.370000  0.085000  8.540000 0.545000 ;
      RECT 8.710000  0.255000  9.040000 0.735000 ;
      RECT 8.790000  1.835000  8.960000 2.635000 ;
      RECT 9.130000  1.665000  9.460000 2.465000 ;
      RECT 9.210000  0.085000  9.470000 0.545000 ;
      RECT 9.630000  1.495000 10.035000 2.635000 ;
      RECT 9.645000  0.255000 10.035000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__o32ai_4
MACRO sky130_fd_sc_hd__lpflow_inputisolatch_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputisolatch_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.750000 0.765000 2.125000 1.095000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.690000 0.415000 4.975000 0.745000 ;
        RECT 4.690000 1.670000 4.975000 2.455000 ;
        RECT 4.805000 0.745000 4.975000 1.670000 ;
    END
  END Q
  PIN SLEEP_B
    ANTENNAGATEAREA  0.145500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
    END
  END SLEEP_B
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.130000 ;
      RECT 0.610000  1.130000 0.810000 1.460000 ;
      RECT 0.610000  1.460000 0.780000 1.795000 ;
      RECT 0.980000  0.740000 1.185000 0.910000 ;
      RECT 0.980000  0.910000 1.150000 1.825000 ;
      RECT 0.980000  1.825000 1.185000 1.915000 ;
      RECT 0.980000  1.915000 2.845000 1.965000 ;
      RECT 1.015000  0.345000 1.185000 0.740000 ;
      RECT 1.015000  1.965000 2.845000 2.085000 ;
      RECT 1.015000  2.085000 1.185000 2.465000 ;
      RECT 1.320000  1.240000 1.490000 1.525000 ;
      RECT 1.320000  1.525000 2.335000 1.695000 ;
      RECT 1.455000  0.085000 1.785000 0.465000 ;
      RECT 1.455000  2.255000 1.850000 2.635000 ;
      RECT 2.050000  1.355000 2.335000 1.525000 ;
      RECT 2.295000  0.705000 2.675000 1.035000 ;
      RECT 2.310000  2.255000 3.185000 2.425000 ;
      RECT 2.380000  0.365000 3.040000 0.535000 ;
      RECT 2.505000  1.035000 2.675000 1.575000 ;
      RECT 2.505000  1.575000 2.845000 1.915000 ;
      RECT 2.870000  0.535000 3.040000 0.995000 ;
      RECT 2.870000  0.995000 3.780000 1.165000 ;
      RECT 3.015000  1.165000 3.780000 1.325000 ;
      RECT 3.015000  1.325000 3.185000 2.255000 ;
      RECT 3.265000  0.085000 3.595000 0.530000 ;
      RECT 3.355000  2.135000 3.525000 2.635000 ;
      RECT 3.420000  1.535000 4.125000 1.865000 ;
      RECT 3.835000  0.415000 4.125000 0.745000 ;
      RECT 3.835000  1.865000 4.125000 2.435000 ;
      RECT 3.950000  0.745000 4.125000 1.535000 ;
      RECT 4.295000  0.085000 4.465000 0.715000 ;
      RECT 4.295000  1.570000 4.465000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_inputisolatch_1
MACRO sky130_fd_sc_hd__dlrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.955000 1.765000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.610000 0.345000 5.895000 0.745000 ;
        RECT 5.635000 1.670000 5.895000 2.455000 ;
        RECT 5.725000 0.745000 5.895000 1.670000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.745000 0.345000 4.975000 0.995000 ;
        RECT 4.745000 0.995000 5.075000 1.325000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.325000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  1.795000 0.775000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.170000  0.345000 0.345000 0.635000 ;
      RECT 0.170000  0.635000 0.775000 0.805000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.605000  0.805000 0.775000 1.070000 ;
      RECT 0.605000  1.070000 0.835000 1.400000 ;
      RECT 0.605000  1.400000 0.775000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.235000 2.465000 ;
      RECT 1.430000  1.495000 2.115000 1.665000 ;
      RECT 1.430000  1.665000 1.785000 2.415000 ;
      RECT 1.510000  0.345000 1.705000 0.615000 ;
      RECT 1.510000  0.615000 2.115000 0.765000 ;
      RECT 1.510000  0.765000 2.335000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.945000  0.785000 2.335000 1.095000 ;
      RECT 1.945000  1.095000 2.115000 1.495000 ;
      RECT 1.955000  1.835000 2.245000 2.635000 ;
      RECT 2.445000  1.355000 2.835000 1.625000 ;
      RECT 2.445000  1.625000 2.760000 1.685000 ;
      RECT 2.690000  0.765000 3.245000 1.095000 ;
      RECT 2.810000  2.255000 3.625000 2.425000 ;
      RECT 2.815000  0.365000 3.585000 0.535000 ;
      RECT 2.900000  1.785000 3.265000 1.995000 ;
      RECT 3.005000  1.095000 3.245000 1.635000 ;
      RECT 3.005000  1.635000 3.265000 1.785000 ;
      RECT 3.415000  0.535000 3.585000 0.995000 ;
      RECT 3.415000  0.995000 4.175000 1.165000 ;
      RECT 3.455000  1.165000 4.175000 1.325000 ;
      RECT 3.455000  1.325000 3.625000 2.255000 ;
      RECT 3.755000  0.085000 4.025000 0.610000 ;
      RECT 3.815000  1.535000 5.465000 1.735000 ;
      RECT 3.815000  1.735000 4.965000 1.865000 ;
      RECT 3.930000  2.135000 4.445000 2.635000 ;
      RECT 4.195000  0.295000 4.575000 0.805000 ;
      RECT 4.345000  0.805000 4.575000 1.505000 ;
      RECT 4.345000  1.505000 5.465000 1.535000 ;
      RECT 4.625000  1.865000 4.965000 2.435000 ;
      RECT 5.135000  1.915000 5.465000 2.635000 ;
      RECT 5.155000  0.085000 5.440000 0.715000 ;
      RECT 5.245000  0.995000 5.555000 1.325000 ;
      RECT 5.245000  1.325000 5.465000 1.505000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  1.445000 0.775000 1.615000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  1.785000 1.235000 1.955000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.445000 2.615000 1.615000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.925000  1.785000 3.095000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 0.545000 1.415000 0.835000 1.460000 ;
      RECT 0.545000 1.460000 2.675000 1.600000 ;
      RECT 0.545000 1.600000 0.835000 1.645000 ;
      RECT 1.005000 1.755000 1.295000 1.800000 ;
      RECT 1.005000 1.800000 3.155000 1.940000 ;
      RECT 1.005000 1.940000 1.295000 1.985000 ;
      RECT 2.385000 1.415000 2.675000 1.460000 ;
      RECT 2.385000 1.600000 2.675000 1.645000 ;
      RECT 2.865000 1.755000 3.155000 1.800000 ;
      RECT 2.865000 1.940000 3.155000 1.985000 ;
  END
END sky130_fd_sc_hd__dlrtp_1
MACRO sky130_fd_sc_hd__dlrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.955000 1.795000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.014750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.610000 0.255000 5.965000 0.485000 ;
        RECT 5.680000 1.875000 5.965000 2.465000 ;
        RECT 5.795000 0.485000 5.965000 0.765000 ;
        RECT 5.795000 0.765000 7.275000 1.325000 ;
        RECT 5.795000 1.325000 5.965000 1.875000 ;
        RECT 6.575000 0.255000 6.775000 0.765000 ;
        RECT 6.575000 1.325000 6.775000 2.465000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505000 0.995000 5.145000 1.325000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.360000 2.805000 ;
        RECT 0.515000 2.135000 0.845000 2.635000 ;
        RECT 1.960000 1.835000 2.275000 2.635000 ;
        RECT 3.825000 2.135000 4.115000 2.635000 ;
        RECT 4.305000 2.135000 4.585000 2.635000 ;
        RECT 5.115000 1.875000 5.485000 2.635000 ;
        RECT 6.135000 1.495000 6.405000 2.635000 ;
        RECT 6.945000 1.495000 7.275000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.460000  1.495000 2.145000 1.665000 ;
      RECT 1.460000  1.665000 1.790000 2.415000 ;
      RECT 1.540000  0.345000 1.710000 0.615000 ;
      RECT 1.540000  0.615000 2.145000 0.765000 ;
      RECT 1.540000  0.765000 2.345000 0.785000 ;
      RECT 1.880000  0.085000 2.210000 0.445000 ;
      RECT 1.975000  0.785000 2.345000 1.095000 ;
      RECT 1.975000  1.095000 2.145000 1.495000 ;
      RECT 2.475000  1.355000 2.760000 1.685000 ;
      RECT 2.720000  0.705000 3.100000 1.035000 ;
      RECT 2.845000  0.365000 3.505000 0.535000 ;
      RECT 2.905000  2.255000 3.655000 2.425000 ;
      RECT 2.930000  1.035000 3.100000 1.575000 ;
      RECT 2.930000  1.575000 3.270000 1.995000 ;
      RECT 3.335000  0.535000 3.505000 0.995000 ;
      RECT 3.335000  0.995000 4.235000 1.165000 ;
      RECT 3.485000  1.165000 4.235000 1.325000 ;
      RECT 3.485000  1.325000 3.655000 2.255000 ;
      RECT 3.745000  0.085000 4.075000 0.530000 ;
      RECT 3.825000  1.535000 5.625000 1.705000 ;
      RECT 3.825000  1.705000 4.945000 1.865000 ;
      RECT 4.265000  0.255000 4.595000 0.655000 ;
      RECT 4.265000  0.655000 5.625000 0.825000 ;
      RECT 4.755000  1.865000 4.945000 2.465000 ;
      RECT 5.100000  0.085000 5.440000 0.485000 ;
      RECT 5.455000  0.825000 5.625000 1.535000 ;
      RECT 6.135000  0.085000 6.405000 0.595000 ;
      RECT 6.945000  0.085000 7.275000 0.595000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.475000  1.445000 2.645000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.935000  1.785000 3.105000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 2.705000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 3.165000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.415000 1.415000 2.705000 1.460000 ;
      RECT 2.415000 1.600000 2.705000 1.645000 ;
      RECT 2.875000 1.755000 3.165000 1.800000 ;
      RECT 2.875000 1.940000 3.165000 1.985000 ;
  END
END sky130_fd_sc_hd__dlrtp_4
MACRO sky130_fd_sc_hd__dlrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 0.955000 1.770000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.595000 0.255000 5.925000 0.485000 ;
        RECT 5.655000 1.875000 5.925000 2.465000 ;
        RECT 5.755000 0.485000 5.925000 0.765000 ;
        RECT 5.755000 0.765000 6.355000 0.865000 ;
        RECT 5.755000 1.425000 6.355000 1.500000 ;
        RECT 5.755000 1.500000 5.925000 1.875000 ;
        RECT 5.760000 1.415000 6.355000 1.425000 ;
        RECT 5.765000 1.410000 6.355000 1.415000 ;
        RECT 5.770000 0.865000 6.355000 0.890000 ;
        RECT 5.775000 1.385000 6.355000 1.410000 ;
        RECT 5.785000 0.890000 6.355000 1.385000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.480000 0.995000 4.815000 1.035000 ;
        RECT 4.480000 1.035000 5.240000 1.325000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.435000  1.495000 2.120000 1.665000 ;
      RECT 1.435000  1.665000 1.785000 2.415000 ;
      RECT 1.515000  0.345000 1.705000 0.615000 ;
      RECT 1.515000  0.615000 2.120000 0.765000 ;
      RECT 1.515000  0.765000 2.335000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.950000  0.785000 2.335000 1.095000 ;
      RECT 1.950000  1.095000 2.120000 1.495000 ;
      RECT 1.955000  1.835000 2.250000 2.635000 ;
      RECT 2.450000  1.355000 2.755000 1.685000 ;
      RECT 2.585000  0.735000 3.100000 1.040000 ;
      RECT 2.770000  0.365000 3.445000 0.535000 ;
      RECT 2.770000  2.255000 3.580000 2.425000 ;
      RECT 2.905000  1.780000 3.265000 1.910000 ;
      RECT 2.905000  1.910000 3.175000 1.995000 ;
      RECT 2.930000  1.040000 3.100000 1.570000 ;
      RECT 2.930000  1.570000 3.265000 1.780000 ;
      RECT 3.270000  0.535000 3.445000 0.995000 ;
      RECT 3.270000  0.995000 4.220000 1.325000 ;
      RECT 3.410000  2.000000 3.605000 2.085000 ;
      RECT 3.410000  2.085000 3.580000 2.255000 ;
      RECT 3.415000  1.995000 3.605000 2.000000 ;
      RECT 3.420000  1.985000 3.605000 1.995000 ;
      RECT 3.435000  1.325000 3.605000 1.985000 ;
      RECT 3.720000  0.085000 4.060000 0.530000 ;
      RECT 3.750000  2.175000 4.090000 2.635000 ;
      RECT 3.775000  1.535000 5.585000 1.705000 ;
      RECT 3.775000  1.705000 4.970000 1.865000 ;
      RECT 4.240000  0.255000 4.580000 0.655000 ;
      RECT 4.240000  0.655000 5.095000 0.695000 ;
      RECT 4.240000  0.695000 5.585000 0.825000 ;
      RECT 4.280000  2.135000 4.560000 2.635000 ;
      RECT 4.800000  1.865000 4.970000 2.465000 ;
      RECT 4.955000  0.825000 5.585000 0.865000 ;
      RECT 5.140000  1.875000 5.485000 2.635000 ;
      RECT 5.255000  0.085000 5.425000 0.525000 ;
      RECT 5.415000  0.865000 5.585000 0.995000 ;
      RECT 5.415000  0.995000 5.615000 1.325000 ;
      RECT 5.415000  1.325000 5.585000 1.535000 ;
      RECT 6.095000  0.085000 6.355000 0.595000 ;
      RECT 6.095000  1.670000 6.355000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.450000  1.445000 2.620000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.925000  1.785000 3.095000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 2.680000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 3.155000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.390000 1.415000 2.680000 1.460000 ;
      RECT 2.390000 1.600000 2.680000 1.645000 ;
      RECT 2.865000 1.755000 3.155000 1.800000 ;
      RECT 2.865000 1.940000 3.155000 1.985000 ;
  END
END sky130_fd_sc_hd__dlrtp_2
MACRO sky130_fd_sc_hd__and2_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.185000 0.430000 1.955000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.940000 1.080000 1.270000 1.615000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.280900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.560000 0.255000 2.215000 0.525000 ;
        RECT 1.790000 1.835000 2.215000 2.465000 ;
        RECT 1.950000 0.525000 2.215000 1.835000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.160000  2.175000 0.430000 2.635000 ;
      RECT 0.185000  0.280000 0.490000 0.695000 ;
      RECT 0.185000  0.695000 1.780000 0.910000 ;
      RECT 0.185000  0.910000 0.770000 0.950000 ;
      RECT 0.600000  0.950000 0.770000 2.135000 ;
      RECT 0.600000  2.135000 0.865000 2.465000 ;
      RECT 0.950000  0.085000 1.390000 0.525000 ;
      RECT 1.110000  1.835000 1.620000 2.635000 ;
      RECT 1.450000  0.910000 1.780000 1.435000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__and2_0
MACRO sky130_fd_sc_hd__and2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.775000 1.325000 ;
        RECT 0.085000 1.325000 0.400000 1.765000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.075000 1.335000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.643500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.665000 0.255000 2.215000 0.545000 ;
        RECT 1.765000 1.915000 2.215000 2.465000 ;
        RECT 1.965000 0.545000 2.215000 1.915000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.285000  0.355000 0.615000 0.715000 ;
      RECT 0.285000  0.715000 1.675000 0.905000 ;
      RECT 0.285000  1.965000 0.565000 2.635000 ;
      RECT 0.735000  1.575000 1.675000 1.745000 ;
      RECT 0.735000  1.745000 1.035000 2.295000 ;
      RECT 1.245000  0.085000 1.495000 0.545000 ;
      RECT 1.245000  1.915000 1.575000 2.635000 ;
      RECT 1.505000  0.905000 1.675000 0.995000 ;
      RECT 1.505000  0.995000 1.795000 1.325000 ;
      RECT 1.505000  1.325000 1.675000 1.575000 ;
      RECT 2.385000  0.085000 2.675000 0.885000 ;
      RECT 2.385000  1.495000 2.675000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__and2_2
MACRO sky130_fd_sc_hd__and2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.995000 0.435000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.995000 0.980000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.515000 1.720000 0.615000 ;
        RECT 1.530000 0.615000 3.135000 0.845000 ;
        RECT 1.530000 1.535000 3.135000 1.760000 ;
        RECT 1.530000 1.760000 1.720000 2.465000 ;
        RECT 2.390000 0.255000 2.580000 0.615000 ;
        RECT 2.390000 1.760000 3.135000 1.765000 ;
        RECT 2.390000 1.765000 2.580000 2.465000 ;
        RECT 2.855000 0.845000 3.135000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.095000  0.255000 0.425000 0.615000 ;
      RECT 0.095000  0.615000 1.360000 0.805000 ;
      RECT 0.095000  1.880000 0.425000 2.635000 ;
      RECT 0.605000  1.580000 1.360000 1.750000 ;
      RECT 0.605000  1.750000 0.785000 2.465000 ;
      RECT 0.955000  0.085000 1.285000 0.445000 ;
      RECT 0.990000  1.935000 1.320000 2.635000 ;
      RECT 1.150000  0.805000 1.360000 1.020000 ;
      RECT 1.150000  1.020000 2.685000 1.355000 ;
      RECT 1.150000  1.355000 1.360000 1.580000 ;
      RECT 1.890000  0.085000 2.220000 0.445000 ;
      RECT 1.890000  1.935000 2.220000 2.635000 ;
      RECT 2.750000  0.085000 3.080000 0.445000 ;
      RECT 2.750000  1.935000 3.080000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__and2_4
MACRO sky130_fd_sc_hd__and2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 0.775000 1.325000 ;
        RECT 0.100000 1.325000 0.365000 1.685000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.075000 1.335000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.657000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655000 0.255000 2.215000 0.545000 ;
        RECT 1.755000 1.915000 2.215000 2.465000 ;
        RECT 1.965000 0.545000 2.215000 1.915000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.285000  0.355000 0.615000 0.715000 ;
      RECT 0.285000  0.715000 1.675000 0.905000 ;
      RECT 0.285000  1.965000 0.565000 2.635000 ;
      RECT 0.735000  1.575000 1.675000 1.745000 ;
      RECT 0.735000  1.745000 1.035000 2.295000 ;
      RECT 1.235000  0.085000 1.485000 0.545000 ;
      RECT 1.235000  1.915000 1.565000 2.635000 ;
      RECT 1.505000  0.905000 1.675000 0.995000 ;
      RECT 1.505000  0.995000 1.795000 1.325000 ;
      RECT 1.505000  1.325000 1.675000 1.575000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__and2_1
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.402500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.290000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 2.370000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 6.440000 5.680000 ;
      LAYER pwell ;
        RECT 0.145000 4.595000 0.315000 5.120000 ;
        RECT 5.925000 4.595000 6.095000 5.120000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.500000 6.170000 3.640000 ;
        RECT 0.080000 3.455000 0.370000 3.500000 ;
        RECT 0.080000 3.640000 0.370000 3.685000 ;
        RECT 5.870000 3.455000 6.160000 3.500000 ;
        RECT 5.870000 3.640000 6.160000 3.685000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 4.135000 ;
        RECT  4.250000 1.305000 6.630000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  PIN VPWRIN
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 6.170000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END VPWRIN
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 6.440000 5.525000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  2.985000 0.375000 3.970000 ;
      RECT 0.085000  4.630000 0.375000 5.355000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.290000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.290000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 6.440000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.865000  0.085000 6.155000 0.810000 ;
      RECT 5.865000  2.985000 6.155000 3.955000 ;
      RECT 5.865000  4.630000 6.155000 5.355000 ;
    LAYER mcon ;
      RECT 0.140000  3.485000 0.310000 3.655000 ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 5.930000  3.485000 6.100000 3.655000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 6.440000 0.240000 ;
    LAYER pwell ;
      RECT 0.145000 0.320000 0.315000 0.845000 ;
      RECT 5.925000 0.320000 6.095000 0.845000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.610500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.255000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 2.370000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 6.440000 5.680000 ;
      LAYER pwell ;
        RECT 0.145000 4.595000 0.315000 5.120000 ;
        RECT 6.125000 4.595000 6.295000 5.120000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.500000 6.300000 3.640000 ;
        RECT 0.080000 3.455000 0.370000 3.500000 ;
        RECT 0.080000 3.640000 0.370000 3.685000 ;
        RECT 6.010000 3.455000 6.300000 3.500000 ;
        RECT 6.010000 3.640000 6.300000 3.685000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 4.135000 ;
        RECT  4.250000 1.305000 6.630000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  PIN VPWRIN
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 6.370000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END VPWRIN
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 6.440000 5.525000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  2.985000 0.375000 3.970000 ;
      RECT 0.085000  4.630000 0.375000 5.355000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.255000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.255000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 6.440000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.825000  0.085000 6.155000 0.900000 ;
      RECT 5.905000  1.610000 6.075000 2.635000 ;
      RECT 6.065000  2.985000 6.355000 3.955000 ;
      RECT 6.065000  4.630000 6.355000 5.355000 ;
    LAYER mcon ;
      RECT 0.140000  3.485000 0.310000 3.655000 ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 6.070000  3.485000 6.240000 3.655000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 6.440000 0.240000 ;
    LAYER pwell ;
      RECT 0.145000 0.320000 0.315000 0.845000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.072500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.255000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 1.085000 ;
        RECT 5.360000 1.085000 6.555000 1.410000 ;
        RECT 5.360000 1.410000 5.635000 2.370000 ;
        RECT 6.280000 1.410000 6.555000 2.370000 ;
        RECT 6.335000 0.255000 6.555000 1.085000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 7.360000 5.680000 ;
      LAYER pwell ;
        RECT 0.145000 4.595000 0.315000 5.120000 ;
        RECT 7.045000 4.595000 7.215000 5.120000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.500000 7.290000 3.640000 ;
        RECT 0.080000 3.455000 0.370000 3.500000 ;
        RECT 0.080000 3.640000 0.370000 3.685000 ;
        RECT 6.930000 3.455000 7.220000 3.500000 ;
        RECT 6.930000 3.640000 7.220000 3.685000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 4.135000 ;
        RECT  4.250000 1.305000 7.405000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  PIN VPWRIN
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 7.290000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END VPWRIN
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 7.360000 5.525000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  2.985000 0.375000 3.970000 ;
      RECT 0.085000  4.630000 0.375000 5.355000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.255000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.255000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 7.360000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.825000  0.085000 6.155000 0.845000 ;
      RECT 5.905000  1.610000 6.075000 2.635000 ;
      RECT 6.755000  0.085000 7.005000 0.925000 ;
      RECT 6.755000  1.610000 6.935000 2.635000 ;
      RECT 6.985000  2.985000 7.275000 3.955000 ;
      RECT 6.985000  4.630000 7.275000 5.355000 ;
    LAYER mcon ;
      RECT 0.140000  3.485000 0.310000 3.655000 ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.585000  5.355000 6.755000 5.525000 ;
      RECT 6.990000  3.485000 7.160000 3.655000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.045000  5.355000 7.215000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 7.360000 0.240000 ;
    LAYER pwell ;
      RECT 0.145000 0.320000 0.315000 0.845000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4
MACRO sky130_fd_sc_hd__dlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlclkp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.765000 1.950000 1.015000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.039500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.040000 0.255000 6.460000 0.545000 ;
        RECT 6.040000 1.835000 7.300000 2.005000 ;
        RECT 6.040000 2.005000 6.370000 2.455000 ;
        RECT 6.290000 0.545000 6.460000 0.715000 ;
        RECT 6.290000 0.715000 7.300000 0.885000 ;
        RECT 6.585000 1.785000 7.300000 1.835000 ;
        RECT 6.750000 0.885000 7.300000 1.785000 ;
        RECT 6.970000 0.255000 7.300000 0.715000 ;
        RECT 6.970000 2.005000 7.300000 2.465000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.406500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
      LAYER mcon ;
        RECT 0.150000 1.105000 0.320000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.230000 1.055000 5.740000 1.325000 ;
      LAYER mcon ;
        RECT 5.230000 1.105000 5.400000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.090000 1.075000 0.380000 1.120000 ;
        RECT 0.090000 1.120000 5.460000 1.260000 ;
        RECT 0.090000 1.260000 0.380000 1.305000 ;
        RECT 5.170000 1.075000 5.460000 1.120000 ;
        RECT 5.170000 1.260000 5.460000 1.305000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.780000 0.805000 ;
      RECT 0.085000  1.795000 0.780000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.280000 1.355000 ;
      RECT 1.015000  1.355000 2.335000 1.585000 ;
      RECT 1.015000  1.585000 1.240000 2.465000 ;
      RECT 1.450000  0.085000 1.785000 0.465000 ;
      RECT 1.450000  2.195000 1.815000 2.635000 ;
      RECT 1.525000  1.785000 1.695000 1.855000 ;
      RECT 1.525000  1.855000 2.845000 1.905000 ;
      RECT 1.525000  1.905000 2.735000 2.025000 ;
      RECT 2.045000  1.585000 2.335000 1.685000 ;
      RECT 2.290000  0.705000 2.735000 1.035000 ;
      RECT 2.415000  0.365000 3.075000 0.535000 ;
      RECT 2.475000  2.195000 3.165000 2.425000 ;
      RECT 2.505000  1.575000 2.845000 1.855000 ;
      RECT 2.565000  1.035000 2.735000 1.575000 ;
      RECT 2.905000  0.535000 3.075000 0.995000 ;
      RECT 2.905000  0.995000 3.775000 1.165000 ;
      RECT 2.915000  2.060000 3.185000 2.090000 ;
      RECT 2.915000  2.090000 3.180000 2.105000 ;
      RECT 2.915000  2.105000 3.165000 2.195000 ;
      RECT 2.980000  2.015000 3.185000 2.060000 ;
      RECT 3.015000  1.165000 3.775000 1.325000 ;
      RECT 3.015000  1.325000 3.185000 2.015000 ;
      RECT 3.315000  0.085000 3.650000 0.530000 ;
      RECT 3.335000  2.175000 3.695000 2.635000 ;
      RECT 3.355000  1.535000 4.115000 1.865000 ;
      RECT 3.895000  0.415000 4.115000 0.745000 ;
      RECT 3.895000  1.865000 4.115000 2.435000 ;
      RECT 3.945000  0.745000 4.115000 0.995000 ;
      RECT 3.945000  0.995000 4.720000 1.325000 ;
      RECT 3.945000  1.325000 4.115000 1.535000 ;
      RECT 4.295000  0.085000 4.580000 0.715000 ;
      RECT 4.295000  2.010000 4.580000 2.635000 ;
      RECT 4.750000  0.290000 5.060000 0.715000 ;
      RECT 4.750000  0.715000 6.120000 0.825000 ;
      RECT 4.750000  1.495000 6.140000 1.665000 ;
      RECT 4.750000  1.665000 5.035000 2.465000 ;
      RECT 4.890000  0.825000 6.120000 0.885000 ;
      RECT 4.890000  0.885000 5.060000 1.495000 ;
      RECT 5.575000  1.835000 5.840000 2.635000 ;
      RECT 5.590000  0.085000 5.870000 0.545000 ;
      RECT 5.910000  0.885000 6.120000 1.055000 ;
      RECT 5.910000  1.055000 6.580000 1.290000 ;
      RECT 5.910000  1.290000 6.140000 1.495000 ;
      RECT 6.540000  2.175000 6.800000 2.635000 ;
      RECT 6.630000  0.085000 6.800000 0.545000 ;
      RECT 7.470000  0.085000 7.735000 0.885000 ;
      RECT 7.470000  1.485000 7.735000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.785000 0.780000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.755000 0.840000 1.800000 ;
      RECT 0.550000 1.800000 1.755000 1.940000 ;
      RECT 0.550000 1.940000 0.840000 1.985000 ;
      RECT 1.465000 1.755000 1.755000 1.800000 ;
      RECT 1.465000 1.940000 1.755000 1.985000 ;
  END
END sky130_fd_sc_hd__dlclkp_4
MACRO sky130_fd_sc_hd__dlclkp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlclkp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 1.435000 2.215000 1.685000 ;
        RECT 1.985000 0.285000 2.215000 1.435000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.060000 0.255000 6.360000 0.595000 ;
        RECT 6.095000 1.495000 6.360000 2.455000 ;
        RECT 6.165000 0.595000 6.360000 1.495000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
      LAYER mcon ;
        RECT 0.150000 1.105000 0.320000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.210000 1.105000 5.485000 1.435000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.090000 1.075000 0.380000 1.120000 ;
        RECT 0.090000 1.120000 5.440000 1.260000 ;
        RECT 0.090000 1.260000 0.380000 1.305000 ;
        RECT 5.150000 1.075000 5.440000 1.120000 ;
        RECT 5.150000 1.260000 5.440000 1.305000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 0.995000 1.355000 ;
        RECT -0.190000 1.355000 7.090000 2.910000 ;
        RECT  2.625000 1.305000 7.090000 1.355000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.175000  0.260000 0.345000 0.615000 ;
      RECT 0.175000  0.615000 0.780000 0.785000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.785000 0.780000 1.060000 ;
      RECT 0.610000  1.060000 0.840000 1.390000 ;
      RECT 0.610000  1.390000 0.780000 1.795000 ;
      RECT 1.015000  0.260000 1.280000 1.855000 ;
      RECT 1.015000  1.855000 2.645000 2.025000 ;
      RECT 1.015000  2.025000 1.240000 2.465000 ;
      RECT 1.455000  2.195000 1.820000 2.635000 ;
      RECT 1.485000  0.085000 1.815000 0.905000 ;
      RECT 2.395000  0.815000 3.225000 0.985000 ;
      RECT 2.395000  0.985000 2.645000 1.855000 ;
      RECT 2.480000  2.255000 3.230000 2.425000 ;
      RECT 2.795000  0.390000 3.725000 0.560000 ;
      RECT 3.060000  1.155000 4.180000 1.325000 ;
      RECT 3.060000  1.325000 3.230000 2.255000 ;
      RECT 3.400000  2.135000 3.700000 2.635000 ;
      RECT 3.435000  1.535000 4.735000 1.840000 ;
      RECT 3.435000  1.840000 4.135000 1.865000 ;
      RECT 3.555000  0.560000 3.725000 0.995000 ;
      RECT 3.555000  0.995000 4.180000 1.155000 ;
      RECT 3.895000  0.085000 4.145000 0.610000 ;
      RECT 3.915000  1.865000 4.135000 2.435000 ;
      RECT 4.315000  0.255000 4.585000 0.615000 ;
      RECT 4.315000  2.010000 4.600000 2.635000 ;
      RECT 4.350000  0.615000 4.585000 0.995000 ;
      RECT 4.350000  0.995000 4.735000 1.535000 ;
      RECT 4.835000  0.290000 5.150000 0.620000 ;
      RECT 4.930000  0.620000 5.150000 0.765000 ;
      RECT 4.930000  0.765000 5.995000 0.935000 ;
      RECT 5.010000  1.725000 5.925000 1.895000 ;
      RECT 5.010000  1.895000 5.340000 2.465000 ;
      RECT 5.575000  2.130000 5.925000 2.635000 ;
      RECT 5.675000  0.085000 5.845000 0.545000 ;
      RECT 5.755000  0.935000 5.995000 1.325000 ;
      RECT 5.755000  1.325000 5.925000 1.725000 ;
      RECT 6.530000  0.085000 6.810000 0.885000 ;
      RECT 6.530000  1.485000 6.810000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
END sky130_fd_sc_hd__dlclkp_2
MACRO sky130_fd_sc_hd__dlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.435000 2.185000 1.685000 ;
        RECT 1.985000 0.385000 2.185000 1.435000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055000 0.255000 6.355000 0.595000 ;
        RECT 6.090000 1.495000 6.355000 2.455000 ;
        RECT 6.170000 0.595000 6.355000 1.495000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
      LAYER mcon ;
        RECT 0.145000 1.105000 0.315000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.190000 1.105000 5.510000 1.435000 ;
      LAYER mcon ;
        RECT 5.210000 1.105000 5.380000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085000 1.075000 0.380000 1.120000 ;
        RECT 0.085000 1.120000 5.440000 1.260000 ;
        RECT 0.085000 1.260000 0.380000 1.305000 ;
        RECT 5.150000 1.075000 5.440000 1.120000 ;
        RECT 5.150000 1.260000 5.440000 1.305000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 0.995000 1.355000 ;
        RECT -0.190000 1.355000 6.630000 2.910000 ;
        RECT  2.620000 1.305000 6.630000 1.355000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.260000 0.345000 0.615000 ;
      RECT 0.175000  0.615000 0.780000 0.785000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.785000 0.780000 1.060000 ;
      RECT 0.610000  1.060000 0.840000 1.390000 ;
      RECT 0.610000  1.390000 0.780000 1.795000 ;
      RECT 1.015000  0.260000 1.280000 1.855000 ;
      RECT 1.015000  1.855000 2.590000 2.025000 ;
      RECT 1.015000  2.025000 1.240000 2.465000 ;
      RECT 1.450000  2.195000 1.815000 2.635000 ;
      RECT 1.480000  0.085000 1.810000 0.905000 ;
      RECT 2.390000  0.815000 3.220000 0.985000 ;
      RECT 2.390000  0.985000 2.590000 1.855000 ;
      RECT 2.475000  2.255000 3.225000 2.425000 ;
      RECT 2.790000  0.390000 3.725000 0.560000 ;
      RECT 3.055000  1.155000 4.175000 1.325000 ;
      RECT 3.055000  1.325000 3.225000 2.255000 ;
      RECT 3.395000  2.135000 3.695000 2.635000 ;
      RECT 3.430000  1.535000 4.710000 1.840000 ;
      RECT 3.430000  1.840000 4.130000 1.865000 ;
      RECT 3.555000  0.560000 3.725000 0.995000 ;
      RECT 3.555000  0.995000 4.175000 1.155000 ;
      RECT 3.895000  0.085000 4.145000 0.610000 ;
      RECT 3.910000  1.865000 4.130000 2.435000 ;
      RECT 4.310000  2.010000 4.595000 2.635000 ;
      RECT 4.320000  0.255000 4.580000 0.615000 ;
      RECT 4.345000  0.615000 4.580000 0.995000 ;
      RECT 4.345000  0.995000 4.740000 1.325000 ;
      RECT 4.345000  1.325000 4.710000 1.535000 ;
      RECT 4.840000  0.290000 5.155000 0.620000 ;
      RECT 4.935000  0.620000 5.155000 0.765000 ;
      RECT 4.935000  0.765000 6.000000 0.935000 ;
      RECT 5.005000  1.725000 5.920000 1.895000 ;
      RECT 5.005000  1.895000 5.335000 2.465000 ;
      RECT 5.570000  2.130000 5.920000 2.635000 ;
      RECT 5.670000  0.085000 5.840000 0.545000 ;
      RECT 5.750000  0.935000 6.000000 1.325000 ;
      RECT 5.750000  1.325000 5.920000 1.725000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__dlclkp_1
MACRO sky130_fd_sc_hd__or4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.490000 0.995000 1.895000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 2.125000 1.745000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 0.995000 1.320000 1.615000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.755000 0.440000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 0.415000 2.675000 0.760000 ;
        RECT 2.405000 1.495000 2.675000 2.465000 ;
        RECT 2.505000 0.760000 2.675000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  1.495000 0.410000 1.785000 ;
      RECT 0.090000  1.785000 1.680000 1.955000 ;
      RECT 0.095000  0.085000 0.425000 0.585000 ;
      RECT 0.625000  0.305000 0.795000 0.655000 ;
      RECT 0.625000  0.655000 2.235000 0.825000 ;
      RECT 0.995000  0.085000 1.325000 0.485000 ;
      RECT 1.495000  0.305000 1.665000 0.655000 ;
      RECT 1.510000  1.495000 2.235000 1.665000 ;
      RECT 1.510000  1.665000 1.680000 1.785000 ;
      RECT 1.835000  0.085000 2.215000 0.485000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
      RECT 2.065000  0.825000 2.235000 0.995000 ;
      RECT 2.065000  0.995000 2.335000 1.325000 ;
      RECT 2.065000  1.325000 2.235000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__or4_1
MACRO sky130_fd_sc_hd__or4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.840000 0.995000 2.010000 1.445000 ;
        RECT 1.840000 1.445000 2.275000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.280000 0.995000 1.610000 1.450000 ;
        RECT 1.400000 1.450000 1.610000 1.785000 ;
        RECT 1.400000 1.785000 1.720000 2.375000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.880000 0.995000 1.050000 1.620000 ;
        RECT 0.880000 1.620000 1.230000 2.375000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.755000 0.370000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.480000 1.455000 4.055000 1.625000 ;
        RECT 2.480000 1.625000 2.730000 2.465000 ;
        RECT 2.520000 0.255000 2.770000 0.725000 ;
        RECT 2.520000 0.725000 4.055000 0.905000 ;
        RECT 3.280000 0.255000 3.610000 0.725000 ;
        RECT 3.320000 1.625000 3.570000 2.465000 ;
        RECT 3.810000 0.905000 4.055000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.115000  1.495000 0.710000 1.665000 ;
      RECT 0.115000  1.665000 0.450000 2.450000 ;
      RECT 0.120000  0.085000 0.370000 0.585000 ;
      RECT 0.540000  0.655000 2.350000 0.825000 ;
      RECT 0.540000  0.825000 0.710000 1.495000 ;
      RECT 0.700000  0.305000 0.870000 0.655000 ;
      RECT 1.070000  0.085000 1.400000 0.485000 ;
      RECT 1.570000  0.305000 1.740000 0.655000 ;
      RECT 1.960000  0.085000 2.340000 0.485000 ;
      RECT 2.005000  1.795000 2.255000 2.635000 ;
      RECT 2.180000  0.825000 2.350000 1.075000 ;
      RECT 2.180000  1.075000 3.640000 1.245000 ;
      RECT 2.900000  1.795000 3.150000 2.635000 ;
      RECT 2.940000  0.085000 3.110000 0.555000 ;
      RECT 3.740000  1.795000 3.990000 2.635000 ;
      RECT 3.780000  0.085000 3.950000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__or4_4
MACRO sky130_fd_sc_hd__or4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.490000 0.995000 1.895000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 2.125000 1.745000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 0.995000 1.320000 1.615000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.755000 0.440000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 0.415000 2.680000 0.760000 ;
        RECT 2.405000 1.495000 2.680000 2.465000 ;
        RECT 2.510000 0.760000 2.680000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.495000 0.410000 1.785000 ;
      RECT 0.085000  1.785000 1.680000 1.955000 ;
      RECT 0.090000  0.085000 0.425000 0.585000 ;
      RECT 0.625000  0.305000 0.795000 0.655000 ;
      RECT 0.625000  0.655000 2.235000 0.825000 ;
      RECT 0.995000  0.085000 1.325000 0.485000 ;
      RECT 1.495000  0.305000 1.665000 0.655000 ;
      RECT 1.510000  1.495000 2.235000 1.665000 ;
      RECT 1.510000  1.665000 1.680000 1.785000 ;
      RECT 1.835000  0.085000 2.215000 0.485000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
      RECT 2.065000  0.825000 2.235000 0.995000 ;
      RECT 2.065000  0.995000 2.340000 1.325000 ;
      RECT 2.065000  1.325000 2.235000 1.495000 ;
      RECT 2.850000  0.085000 3.020000 1.000000 ;
      RECT 2.850000  1.455000 3.020000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__or4_2
MACRO sky130_fd_sc_hd__dlxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.470250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.150000 0.415000 5.435000 0.745000 ;
        RECT 5.150000 1.670000 5.435000 2.455000 ;
        RECT 5.265000 0.745000 5.435000 1.670000 ;
    END
  END Q
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 1.685000 ;
      RECT 2.715000  0.705000 3.095000 1.035000 ;
      RECT 2.770000  2.255000 3.605000 2.425000 ;
      RECT 2.840000  0.365000 3.500000 0.535000 ;
      RECT 2.925000  1.035000 3.095000 1.575000 ;
      RECT 2.925000  1.575000 3.265000 1.995000 ;
      RECT 3.330000  0.535000 3.500000 0.995000 ;
      RECT 3.330000  0.995000 4.175000 1.165000 ;
      RECT 3.435000  1.165000 4.175000 1.325000 ;
      RECT 3.435000  1.325000 3.605000 2.255000 ;
      RECT 3.685000  0.085000 4.015000 0.530000 ;
      RECT 3.775000  2.135000 3.945000 2.635000 ;
      RECT 3.840000  1.535000 4.515000 1.865000 ;
      RECT 4.295000  0.415000 4.515000 0.745000 ;
      RECT 4.295000  1.865000 4.515000 2.435000 ;
      RECT 4.345000  0.745000 4.515000 0.995000 ;
      RECT 4.345000  0.995000 5.095000 1.325000 ;
      RECT 4.345000  1.325000 4.515000 1.535000 ;
      RECT 4.695000  0.085000 4.900000 0.715000 ;
      RECT 4.695000  1.570000 4.900000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.445000 2.640000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.785000 3.100000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 2.700000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 3.160000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.415000 2.700000 1.460000 ;
      RECT 2.410000 1.600000 2.700000 1.645000 ;
      RECT 2.870000 1.755000 3.160000 1.800000 ;
      RECT 2.870000 1.940000 3.160000 1.985000 ;
  END
END sky130_fd_sc_hd__dlxtp_1
MACRO sky130_fd_sc_hd__and4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.450000 1.675000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 0.420000 1.800000 1.695000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 0.420000 2.295000 1.695000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485000 0.665000 2.825000 1.695000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.255000 0.295000 3.590000 0.340000 ;
        RECT 3.255000 0.340000 3.595000 0.805000 ;
        RECT 3.335000 1.495000 3.595000 2.465000 ;
        RECT 3.425000 0.805000 3.595000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.170000  0.255000 0.345000 0.655000 ;
      RECT 0.170000  0.655000 0.800000 0.825000 ;
      RECT 0.170000  1.845000 0.800000 2.015000 ;
      RECT 0.170000  2.015000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.195000 0.845000 2.635000 ;
      RECT 0.630000  0.825000 0.800000 0.995000 ;
      RECT 0.630000  0.995000 0.980000 1.325000 ;
      RECT 0.630000  1.325000 0.800000 1.845000 ;
      RECT 1.090000  0.255000 1.320000 0.585000 ;
      RECT 1.150000  0.585000 1.320000 1.875000 ;
      RECT 1.150000  1.875000 3.165000 2.045000 ;
      RECT 1.150000  2.045000 1.320000 2.465000 ;
      RECT 1.555000  2.225000 2.225000 2.635000 ;
      RECT 2.440000  2.045000 2.610000 2.465000 ;
      RECT 2.755000  0.085000 3.085000 0.465000 ;
      RECT 2.810000  2.225000 3.140000 2.635000 ;
      RECT 2.995000  0.995000 3.255000 1.325000 ;
      RECT 2.995000  1.325000 3.165000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__and4b_1
MACRO sky130_fd_sc_hd__and4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 0.765000 0.790000 1.635000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 0.735000 4.145000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.345000 0.755000 3.555000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 0.995000 3.085000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.980000 0.650000 2.080000 0.820000 ;
        RECT 0.980000 0.820000 1.260000 1.545000 ;
        RECT 0.980000 1.545000 2.160000 1.715000 ;
        RECT 1.070000 0.255000 1.240000 0.650000 ;
        RECT 1.910000 0.255000 2.080000 0.650000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.260000 1.915000 ;
      RECT 0.085000  1.915000 4.900000 2.085000 ;
      RECT 0.085000  2.085000 0.345000 2.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 0.570000  0.085000 0.900000 0.470000 ;
      RECT 1.410000  0.085000 1.740000 0.470000 ;
      RECT 1.410000  2.255000 1.740000 2.635000 ;
      RECT 1.440000  1.075000 2.550000 1.245000 ;
      RECT 2.250000  2.255000 2.580000 2.635000 ;
      RECT 2.285000  0.085000 2.615000 0.445000 ;
      RECT 2.380000  0.615000 2.965000 0.785000 ;
      RECT 2.380000  0.785000 2.550000 1.075000 ;
      RECT 2.380000  1.245000 2.550000 1.545000 ;
      RECT 2.380000  1.545000 4.545000 1.715000 ;
      RECT 2.795000  0.300000 4.965000 0.470000 ;
      RECT 2.795000  0.470000 2.965000 0.615000 ;
      RECT 3.475000  2.255000 3.805000 2.635000 ;
      RECT 4.390000  0.470000 4.965000 0.810000 ;
      RECT 4.635000  2.255000 4.965000 2.635000 ;
      RECT 4.730000  0.995000 4.900000 1.915000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__and4b_4
MACRO sky130_fd_sc_hd__and4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.740000 0.335000 1.630000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.420000 1.745000 1.745000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 0.420000 2.275000 1.695000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.645000 2.775000 1.615000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.503250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.260000 0.255000 3.545000 0.640000 ;
        RECT 3.260000 0.640000 4.055000 0.825000 ;
        RECT 3.340000 1.535000 4.055000 1.745000 ;
        RECT 3.340000 1.745000 3.545000 2.465000 ;
        RECT 3.425000 0.825000 4.055000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.175000  1.830000 0.805000 2.000000 ;
      RECT 0.175000  2.000000 0.345000 2.465000 ;
      RECT 0.515000  2.195000 0.845000 2.635000 ;
      RECT 0.595000  0.255000 0.805000 0.585000 ;
      RECT 0.635000  0.585000 0.805000 0.995000 ;
      RECT 0.635000  0.995000 0.975000 1.325000 ;
      RECT 0.635000  1.325000 0.805000 1.830000 ;
      RECT 1.015000  1.660000 1.315000 1.915000 ;
      RECT 1.015000  1.915000 3.165000 1.965000 ;
      RECT 1.015000  1.965000 2.610000 2.085000 ;
      RECT 1.015000  2.085000 1.185000 2.465000 ;
      RECT 1.095000  0.255000 1.315000 0.585000 ;
      RECT 1.145000  0.585000 1.315000 1.660000 ;
      RECT 1.555000  2.255000 2.225000 2.635000 ;
      RECT 2.440000  1.795000 3.165000 1.915000 ;
      RECT 2.440000  2.085000 2.610000 2.465000 ;
      RECT 2.760000  0.085000 3.090000 0.465000 ;
      RECT 2.840000  2.195000 3.170000 2.635000 ;
      RECT 2.995000  0.995000 3.255000 1.325000 ;
      RECT 2.995000  1.325000 3.165000 1.795000 ;
      RECT 3.715000  0.085000 4.050000 0.465000 ;
      RECT 3.715000  1.915000 4.050000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__and4b_2
MACRO sky130_fd_sc_hd__clkinvlp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinvlp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.330000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.745000 0.425000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.714000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.255000 1.215000 0.680000 ;
        RECT 0.595000 0.680000 0.955000 1.015000 ;
        RECT 0.595000 1.015000 2.015000 1.295000 ;
        RECT 0.595000 1.295000 0.955000 2.465000 ;
        RECT 1.685000 1.295000 2.015000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.575000 ;
      RECT 0.095000  1.495000 0.425000 2.635000 ;
      RECT 1.155000  1.465000 1.485000 2.635000 ;
      RECT 1.675000  0.085000 2.005000 0.775000 ;
      RECT 2.215000  1.465000 2.545000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinvlp_4
MACRO sky130_fd_sc_hd__clkinvlp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinvlp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.995000 0.600000 1.665000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.436750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.810000 0.315000 1.445000 0.750000 ;
        RECT 0.810000 0.750000 1.235000 2.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.225000  1.835000 0.555000 2.625000 ;
      RECT 0.225000  2.625000 1.740000 2.635000 ;
      RECT 0.295000  0.085000 0.625000 0.745000 ;
      RECT 1.440000  1.455000 1.740000 2.625000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinvlp_2
MACRO sky130_fd_sc_hd__sdfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfstp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.88000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.519750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.035000 0.255000 12.365000 0.825000 ;
        RECT 12.035000 1.495000 12.365000 2.450000 ;
        RECT 12.145000 0.825000 12.365000 1.495000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.765000 0.820000 1.675000 ;
      LAYER mcon ;
        RECT 0.605000 1.105000 0.775000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.370000 1.075000 2.700000 1.600000 ;
      LAYER mcon ;
        RECT 2.445000 1.105000 2.615000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545000 1.075000 0.835000 1.120000 ;
        RECT 0.545000 1.120000 2.675000 1.260000 ;
        RECT 0.545000 1.260000 0.835000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.065000 1.765000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.880000 1.425000 9.135000 1.545000 ;
        RECT 8.880000 1.545000 9.945000 1.725000 ;
      LAYER mcon ;
        RECT 8.940000 1.445000 9.110000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.170000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.880000 1.415000 9.170000 1.460000 ;
        RECT 8.880000 1.600000 9.170000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.615000 ;
        RECT 2.905000 1.615000 3.085000 1.960000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 13.070000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.880000 0.085000 ;
      RECT  0.000000  2.635000 12.880000 2.805000 ;
      RECT  0.085000  0.085000  0.700000 0.595000 ;
      RECT  0.085000  1.845000  1.125000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.785000 2.635000 ;
      RECT  0.870000  0.255000  1.625000 0.555000 ;
      RECT  0.870000  0.555000  1.640000 0.575000 ;
      RECT  0.870000  0.575000  1.650000 0.595000 ;
      RECT  0.955000  2.025000  1.125000 2.255000 ;
      RECT  0.955000  2.255000  2.045000 2.465000 ;
      RECT  1.295000  1.845000  1.695000 2.085000 ;
      RECT  1.380000  0.595000  1.660000 0.600000 ;
      RECT  1.395000  0.600000  1.660000 0.605000 ;
      RECT  1.405000  0.605000  1.660000 0.610000 ;
      RECT  1.420000  0.610000  1.660000 0.615000 ;
      RECT  1.430000  0.615000  1.660000 0.620000 ;
      RECT  1.440000  0.620000  1.665000 0.630000 ;
      RECT  1.445000  0.630000  1.665000 0.635000 ;
      RECT  1.460000  0.635000  1.665000 0.645000 ;
      RECT  1.475000  0.645000  1.670000 0.660000 ;
      RECT  1.475000  0.660000  1.675000 0.665000 ;
      RECT  1.495000  0.665000  1.675000 0.705000 ;
      RECT  1.505000  0.705000  1.675000 0.710000 ;
      RECT  1.505000  0.710000  1.695000 1.845000 ;
      RECT  1.825000  0.085000  2.090000 0.545000 ;
      RECT  1.865000  0.715000  2.520000 0.905000 ;
      RECT  1.865000  0.905000  2.200000 1.770000 ;
      RECT  1.865000  1.770000  2.520000 2.085000 ;
      RECT  2.260000  0.255000  2.520000 0.715000 ;
      RECT  2.270000  2.085000  2.520000 2.465000 ;
      RECT  2.690000  0.085000  3.100000 0.555000 ;
      RECT  2.690000  2.140000  2.985000 2.635000 ;
      RECT  3.255000  1.830000  3.995000 1.990000 ;
      RECT  3.255000  1.990000  3.985000 2.000000 ;
      RECT  3.255000  2.000000  3.425000 2.325000 ;
      RECT  3.270000  0.255000  3.455000 0.715000 ;
      RECT  3.270000  0.715000  3.995000 0.885000 ;
      RECT  3.595000  2.275000  3.925000 2.635000 ;
      RECT  3.625000  0.085000  3.955000 0.545000 ;
      RECT  3.735000  0.885000  3.995000 1.830000 ;
      RECT  4.095000  2.135000  4.440000 2.465000 ;
      RECT  4.125000  0.255000  4.335000 0.585000 ;
      RECT  4.165000  0.585000  4.335000 1.090000 ;
      RECT  4.165000  1.090000  4.490000 1.420000 ;
      RECT  4.165000  1.420000  4.440000 2.135000 ;
      RECT  4.505000  0.255000  4.830000 0.920000 ;
      RECT  4.615000  1.590000  4.915000 1.615000 ;
      RECT  4.615000  1.615000  4.830000 2.465000 ;
      RECT  4.660000  0.920000  4.830000 1.445000 ;
      RECT  4.660000  1.445000  4.915000 1.590000 ;
      RECT  5.000000  0.255000  5.440000 1.225000 ;
      RECT  5.000000  1.225000  7.715000 1.275000 ;
      RECT  5.035000  2.135000  5.755000 2.465000 ;
      RECT  5.085000  1.275000  6.475000 1.395000 ;
      RECT  5.205000  1.575000  5.415000 1.955000 ;
      RECT  5.585000  1.395000  5.755000 2.135000 ;
      RECT  5.610000  0.085000  6.095000 0.465000 ;
      RECT  5.645000  0.635000  6.535000 0.805000 ;
      RECT  5.645000  0.805000  5.975000 1.015000 ;
      RECT  5.925000  1.575000  6.095000 1.935000 ;
      RECT  5.925000  1.935000  6.820000 2.105000 ;
      RECT  5.945000  2.275000  6.330000 2.635000 ;
      RECT  6.285000  0.255000  6.535000 0.635000 ;
      RECT  6.305000  0.975000  7.715000 1.225000 ;
      RECT  6.605000  2.105000  6.820000 2.450000 ;
      RECT  6.705000  0.085000  7.715000 0.805000 ;
      RECT  7.060000  2.125000  8.015000 2.635000 ;
      RECT  7.235000  1.670000  8.135000 1.955000 ;
      RECT  7.355000  1.275000  7.715000 1.325000 ;
      RECT  7.885000  0.720000  9.105000 0.905000 ;
      RECT  7.885000  0.905000  8.135000 1.670000 ;
      RECT  8.185000  2.125000  8.990000 2.460000 ;
      RECT  8.425000  1.075000  8.650000 1.905000 ;
      RECT  8.465000  0.275000  9.910000 0.545000 ;
      RECT  8.820000  0.905000  9.105000 1.255000 ;
      RECT  8.820000  1.895000 10.485000 2.065000 ;
      RECT  8.820000  2.065000  8.990000 2.125000 ;
      RECT  9.160000  2.235000  9.490000 2.635000 ;
      RECT  9.320000  0.855000  9.530000 1.195000 ;
      RECT  9.320000  1.195000 10.915000 1.365000 ;
      RECT  9.660000  2.065000  9.965000 2.450000 ;
      RECT  9.710000  0.545000  9.910000 0.785000 ;
      RECT  9.710000  0.785000 10.515000 1.015000 ;
      RECT 10.115000  0.085000 10.365000 0.545000 ;
      RECT 10.155000  1.605000 10.485000 1.895000 ;
      RECT 10.155000  2.235000 10.485000 2.635000 ;
      RECT 10.575000  0.255000 10.915000 0.585000 ;
      RECT 10.655000  1.365000 10.915000 2.465000 ;
      RECT 10.685000  0.585000 10.915000 1.195000 ;
      RECT 11.085000  0.255000 11.345000 0.995000 ;
      RECT 11.085000  0.995000 11.975000 1.325000 ;
      RECT 11.085000  1.325000 11.345000 2.465000 ;
      RECT 11.570000  0.085000 11.865000 0.825000 ;
      RECT 11.570000  1.790000 11.820000 2.635000 ;
      RECT 12.535000  0.085000 12.795000 0.885000 ;
      RECT 12.535000  1.495000 12.795000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.445000  1.695000 1.615000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  1.785000  3.995000 1.955000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.445000  4.915000 1.615000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.560000  1.785000  7.730000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.480000  1.105000  8.650000 1.275000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.975000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.790000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.710000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.685000 1.415000 4.975000 1.460000 ;
      RECT 4.685000 1.600000 4.975000 1.645000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 7.500000 1.755000 7.790000 1.800000 ;
      RECT 7.500000 1.940000 7.790000 1.985000 ;
      RECT 8.420000 1.075000 8.710000 1.120000 ;
      RECT 8.420000 1.260000 8.710000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfstp_2
MACRO sky130_fd_sc_hd__sdfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.42000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995000 0.275000 12.335000 0.825000 ;
        RECT 11.995000 1.495000 12.335000 2.450000 ;
        RECT 12.145000 0.825000 12.335000 1.495000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.765000 0.820000 1.675000 ;
      LAYER mcon ;
        RECT 0.605000 1.105000 0.775000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.370000 1.075000 2.700000 1.600000 ;
      LAYER mcon ;
        RECT 2.445000 1.105000 2.615000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545000 1.075000 0.835000 1.120000 ;
        RECT 0.545000 1.120000 2.675000 1.260000 ;
        RECT 0.545000 1.260000 0.835000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.065000 1.765000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.880000 1.425000 9.135000 1.545000 ;
        RECT 8.880000 1.545000 9.945000 1.725000 ;
      LAYER mcon ;
        RECT 8.940000 1.445000 9.110000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.170000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.880000 1.415000 9.170000 1.460000 ;
        RECT 8.880000 1.600000 9.170000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.615000 ;
        RECT 2.905000 1.615000 3.085000 1.960000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.610000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.085000  0.085000  0.700000 0.595000 ;
      RECT  0.085000  1.845000  1.125000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.785000 2.635000 ;
      RECT  0.870000  0.255000  1.625000 0.555000 ;
      RECT  0.870000  0.555000  1.640000 0.575000 ;
      RECT  0.870000  0.575000  1.650000 0.595000 ;
      RECT  0.955000  2.025000  1.125000 2.255000 ;
      RECT  0.955000  2.255000  2.045000 2.465000 ;
      RECT  1.295000  1.845000  1.695000 2.085000 ;
      RECT  1.380000  0.595000  1.660000 0.600000 ;
      RECT  1.395000  0.600000  1.660000 0.605000 ;
      RECT  1.405000  0.605000  1.660000 0.610000 ;
      RECT  1.420000  0.610000  1.660000 0.615000 ;
      RECT  1.430000  0.615000  1.660000 0.620000 ;
      RECT  1.440000  0.620000  1.665000 0.630000 ;
      RECT  1.445000  0.630000  1.665000 0.635000 ;
      RECT  1.460000  0.635000  1.665000 0.645000 ;
      RECT  1.475000  0.645000  1.670000 0.660000 ;
      RECT  1.475000  0.660000  1.675000 0.665000 ;
      RECT  1.495000  0.665000  1.675000 0.705000 ;
      RECT  1.505000  0.705000  1.675000 0.710000 ;
      RECT  1.505000  0.710000  1.695000 1.845000 ;
      RECT  1.825000  0.085000  2.090000 0.545000 ;
      RECT  1.865000  0.715000  2.520000 0.905000 ;
      RECT  1.865000  0.905000  2.200000 1.770000 ;
      RECT  1.865000  1.770000  2.520000 2.085000 ;
      RECT  2.260000  0.255000  2.520000 0.715000 ;
      RECT  2.270000  2.085000  2.520000 2.465000 ;
      RECT  2.690000  0.085000  3.100000 0.555000 ;
      RECT  2.690000  2.140000  2.985000 2.635000 ;
      RECT  3.255000  1.830000  3.995000 1.990000 ;
      RECT  3.255000  1.990000  3.985000 2.000000 ;
      RECT  3.255000  2.000000  3.425000 2.325000 ;
      RECT  3.270000  0.255000  3.455000 0.715000 ;
      RECT  3.270000  0.715000  3.995000 0.885000 ;
      RECT  3.595000  2.275000  3.925000 2.635000 ;
      RECT  3.625000  0.085000  3.955000 0.545000 ;
      RECT  3.735000  0.885000  3.995000 1.830000 ;
      RECT  4.095000  2.135000  4.440000 2.465000 ;
      RECT  4.125000  0.255000  4.335000 0.585000 ;
      RECT  4.165000  0.585000  4.335000 1.090000 ;
      RECT  4.165000  1.090000  4.490000 1.420000 ;
      RECT  4.165000  1.420000  4.440000 2.135000 ;
      RECT  4.505000  0.255000  4.830000 0.920000 ;
      RECT  4.615000  1.590000  4.915000 1.615000 ;
      RECT  4.615000  1.615000  4.830000 2.465000 ;
      RECT  4.660000  0.920000  4.830000 1.445000 ;
      RECT  4.660000  1.445000  4.915000 1.590000 ;
      RECT  5.000000  0.255000  5.440000 1.225000 ;
      RECT  5.000000  1.225000  7.715000 1.275000 ;
      RECT  5.035000  2.135000  5.755000 2.465000 ;
      RECT  5.085000  1.275000  6.475000 1.395000 ;
      RECT  5.205000  1.575000  5.415000 1.955000 ;
      RECT  5.585000  1.395000  5.755000 2.135000 ;
      RECT  5.610000  0.085000  6.095000 0.465000 ;
      RECT  5.645000  0.635000  6.535000 0.805000 ;
      RECT  5.645000  0.805000  5.975000 1.015000 ;
      RECT  5.925000  1.575000  6.095000 1.935000 ;
      RECT  5.925000  1.935000  6.820000 2.105000 ;
      RECT  5.945000  2.275000  6.330000 2.635000 ;
      RECT  6.285000  0.255000  6.535000 0.635000 ;
      RECT  6.305000  0.975000  7.715000 1.225000 ;
      RECT  6.605000  2.105000  6.820000 2.450000 ;
      RECT  6.705000  0.085000  7.715000 0.805000 ;
      RECT  7.060000  2.125000  8.015000 2.635000 ;
      RECT  7.235000  1.670000  8.135000 1.955000 ;
      RECT  7.355000  1.275000  7.715000 1.325000 ;
      RECT  7.885000  0.720000  9.105000 0.905000 ;
      RECT  7.885000  0.905000  8.135000 1.670000 ;
      RECT  8.185000  2.125000  8.990000 2.460000 ;
      RECT  8.425000  1.075000  8.650000 1.905000 ;
      RECT  8.465000  0.275000  9.910000 0.545000 ;
      RECT  8.820000  0.905000  9.105000 1.255000 ;
      RECT  8.820000  1.895000 10.485000 2.065000 ;
      RECT  8.820000  2.065000  8.990000 2.125000 ;
      RECT  9.160000  2.235000  9.490000 2.635000 ;
      RECT  9.320000  0.855000  9.530000 1.195000 ;
      RECT  9.320000  1.195000 10.915000 1.365000 ;
      RECT  9.660000  2.065000  9.965000 2.450000 ;
      RECT  9.710000  0.545000  9.910000 0.785000 ;
      RECT  9.710000  0.785000 10.515000 1.015000 ;
      RECT 10.115000  0.085000 10.365000 0.545000 ;
      RECT 10.155000  1.605000 10.485000 1.895000 ;
      RECT 10.155000  2.235000 10.485000 2.635000 ;
      RECT 10.575000  0.255000 10.915000 0.585000 ;
      RECT 10.655000  1.365000 10.915000 2.465000 ;
      RECT 10.685000  0.585000 10.915000 1.195000 ;
      RECT 11.085000  0.255000 11.345000 0.995000 ;
      RECT 11.085000  0.995000 11.975000 1.325000 ;
      RECT 11.085000  1.325000 11.345000 2.465000 ;
      RECT 11.515000  0.085000 11.825000 0.825000 ;
      RECT 11.515000  1.790000 11.825000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.445000  1.695000 1.615000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  1.785000  3.995000 1.955000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.445000  4.915000 1.615000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.560000  1.785000  7.730000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.480000  1.105000  8.650000 1.275000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.975000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.790000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.710000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.685000 1.415000 4.975000 1.460000 ;
      RECT 4.685000 1.600000 4.975000 1.645000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 7.500000 1.755000 7.790000 1.800000 ;
      RECT 7.500000 1.940000 7.790000 1.985000 ;
      RECT 8.420000 1.075000 8.710000 1.120000 ;
      RECT 8.420000 1.260000 8.710000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfstp_1
MACRO sky130_fd_sc_hd__sdfstp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfstp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.80000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.040000 0.275000 12.370000 0.825000 ;
        RECT 12.040000 1.495000 12.370000 2.450000 ;
        RECT 12.145000 0.825000 12.370000 1.055000 ;
        RECT 12.145000 1.055000 13.210000 1.325000 ;
        RECT 12.145000 1.325000 12.370000 1.495000 ;
        RECT 12.880000 0.255000 13.210000 1.055000 ;
        RECT 12.880000 1.325000 13.210000 2.465000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.765000 0.820000 1.675000 ;
      LAYER mcon ;
        RECT 0.605000 1.105000 0.775000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.370000 1.075000 2.700000 1.600000 ;
      LAYER mcon ;
        RECT 2.445000 1.105000 2.615000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545000 1.075000 0.835000 1.120000 ;
        RECT 0.545000 1.120000 2.675000 1.260000 ;
        RECT 0.545000 1.260000 0.835000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.065000 1.765000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.880000 1.425000 9.135000 1.545000 ;
        RECT 8.880000 1.545000 9.945000 1.725000 ;
      LAYER mcon ;
        RECT 8.940000 1.445000 9.110000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.170000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.880000 1.415000 9.170000 1.460000 ;
        RECT 8.880000 1.600000 9.170000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.615000 ;
        RECT 2.905000 1.615000 3.085000 1.960000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.800000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 13.990000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.800000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.800000 0.085000 ;
      RECT  0.000000  2.635000 13.800000 2.805000 ;
      RECT  0.085000  0.085000  0.700000 0.595000 ;
      RECT  0.085000  1.845000  1.125000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.785000 2.635000 ;
      RECT  0.870000  0.255000  1.625000 0.555000 ;
      RECT  0.870000  0.555000  1.640000 0.575000 ;
      RECT  0.870000  0.575000  1.650000 0.595000 ;
      RECT  0.955000  2.025000  1.125000 2.255000 ;
      RECT  0.955000  2.255000  2.045000 2.465000 ;
      RECT  1.295000  1.845000  1.695000 2.085000 ;
      RECT  1.380000  0.595000  1.660000 0.600000 ;
      RECT  1.395000  0.600000  1.660000 0.605000 ;
      RECT  1.405000  0.605000  1.660000 0.610000 ;
      RECT  1.420000  0.610000  1.660000 0.615000 ;
      RECT  1.430000  0.615000  1.660000 0.620000 ;
      RECT  1.440000  0.620000  1.665000 0.630000 ;
      RECT  1.445000  0.630000  1.665000 0.635000 ;
      RECT  1.460000  0.635000  1.665000 0.645000 ;
      RECT  1.475000  0.645000  1.670000 0.660000 ;
      RECT  1.475000  0.660000  1.675000 0.665000 ;
      RECT  1.495000  0.665000  1.675000 0.705000 ;
      RECT  1.505000  0.705000  1.675000 0.710000 ;
      RECT  1.505000  0.710000  1.695000 1.845000 ;
      RECT  1.825000  0.085000  2.090000 0.545000 ;
      RECT  1.865000  0.715000  2.520000 0.905000 ;
      RECT  1.865000  0.905000  2.200000 1.770000 ;
      RECT  1.865000  1.770000  2.520000 2.085000 ;
      RECT  2.260000  0.255000  2.520000 0.715000 ;
      RECT  2.270000  2.085000  2.520000 2.465000 ;
      RECT  2.690000  0.085000  3.100000 0.555000 ;
      RECT  2.690000  2.140000  2.985000 2.635000 ;
      RECT  3.255000  1.830000  3.995000 1.990000 ;
      RECT  3.255000  1.990000  3.985000 2.000000 ;
      RECT  3.255000  2.000000  3.425000 2.325000 ;
      RECT  3.270000  0.255000  3.455000 0.715000 ;
      RECT  3.270000  0.715000  3.995000 0.885000 ;
      RECT  3.595000  2.275000  3.925000 2.635000 ;
      RECT  3.625000  0.085000  3.955000 0.545000 ;
      RECT  3.735000  0.885000  3.995000 1.830000 ;
      RECT  4.095000  2.135000  4.440000 2.465000 ;
      RECT  4.125000  0.255000  4.335000 0.585000 ;
      RECT  4.165000  0.585000  4.335000 1.090000 ;
      RECT  4.165000  1.090000  4.490000 1.420000 ;
      RECT  4.165000  1.420000  4.440000 2.135000 ;
      RECT  4.505000  0.255000  4.830000 0.920000 ;
      RECT  4.615000  1.590000  4.915000 1.615000 ;
      RECT  4.615000  1.615000  4.830000 2.465000 ;
      RECT  4.660000  0.920000  4.830000 1.445000 ;
      RECT  4.660000  1.445000  4.915000 1.590000 ;
      RECT  5.000000  0.255000  5.440000 1.225000 ;
      RECT  5.000000  1.225000  7.715000 1.275000 ;
      RECT  5.035000  2.135000  5.755000 2.465000 ;
      RECT  5.085000  1.275000  6.475000 1.395000 ;
      RECT  5.205000  1.575000  5.415000 1.955000 ;
      RECT  5.585000  1.395000  5.755000 2.135000 ;
      RECT  5.610000  0.085000  6.095000 0.465000 ;
      RECT  5.645000  0.635000  6.535000 0.805000 ;
      RECT  5.645000  0.805000  5.975000 1.015000 ;
      RECT  5.925000  1.575000  6.095000 1.935000 ;
      RECT  5.925000  1.935000  6.820000 2.105000 ;
      RECT  5.945000  2.275000  6.330000 2.635000 ;
      RECT  6.285000  0.255000  6.535000 0.635000 ;
      RECT  6.305000  0.975000  7.715000 1.225000 ;
      RECT  6.605000  2.105000  6.820000 2.450000 ;
      RECT  6.705000  0.085000  7.715000 0.805000 ;
      RECT  7.060000  2.125000  8.015000 2.635000 ;
      RECT  7.235000  1.670000  8.135000 1.955000 ;
      RECT  7.355000  1.275000  7.715000 1.325000 ;
      RECT  7.885000  0.720000  9.105000 0.905000 ;
      RECT  7.885000  0.905000  8.135000 1.670000 ;
      RECT  8.185000  2.125000  8.990000 2.460000 ;
      RECT  8.425000  1.075000  8.650000 1.905000 ;
      RECT  8.465000  0.275000  9.910000 0.545000 ;
      RECT  8.820000  0.905000  9.105000 1.255000 ;
      RECT  8.820000  1.895000 10.485000 2.065000 ;
      RECT  8.820000  2.065000  8.990000 2.125000 ;
      RECT  9.160000  2.235000  9.490000 2.635000 ;
      RECT  9.320000  0.855000  9.530000 1.195000 ;
      RECT  9.320000  1.195000 10.915000 1.365000 ;
      RECT  9.660000  2.065000  9.965000 2.450000 ;
      RECT  9.710000  0.545000  9.910000 0.785000 ;
      RECT  9.710000  0.785000 10.515000 1.015000 ;
      RECT 10.115000  0.085000 10.365000 0.545000 ;
      RECT 10.155000  1.605000 10.485000 1.895000 ;
      RECT 10.155000  2.235000 10.485000 2.635000 ;
      RECT 10.575000  0.255000 10.915000 0.585000 ;
      RECT 10.655000  1.365000 10.915000 2.465000 ;
      RECT 10.685000  0.585000 10.915000 1.195000 ;
      RECT 11.085000  0.255000 11.345000 0.995000 ;
      RECT 11.085000  0.995000 11.975000 1.325000 ;
      RECT 11.085000  1.325000 11.345000 2.465000 ;
      RECT 11.515000  0.085000 11.870000 0.825000 ;
      RECT 11.515000  1.495000 11.870000 2.635000 ;
      RECT 12.540000  0.085000 12.710000 0.885000 ;
      RECT 12.540000  1.495000 12.710000 2.635000 ;
      RECT 13.380000  0.085000 13.715000 0.885000 ;
      RECT 13.380000  1.495000 13.715000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.445000  1.695000 1.615000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  1.785000  3.995000 1.955000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.445000  4.915000 1.615000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.560000  1.785000  7.730000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.480000  1.105000  8.650000 1.275000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.975000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.790000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.710000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.685000 1.415000 4.975000 1.460000 ;
      RECT 4.685000 1.600000 4.975000 1.645000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 7.500000 1.755000 7.790000 1.800000 ;
      RECT 7.500000 1.940000 7.790000 1.985000 ;
      RECT 8.420000 1.075000 8.710000 1.120000 ;
      RECT 8.420000 1.260000 8.710000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfstp_4
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.576000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.065000 1.305000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.662600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.460000 1.755000 1.630000 ;
        RECT 0.155000 1.630000 0.375000 2.435000 ;
        RECT 1.025000 0.280000 1.250000 0.725000 ;
        RECT 1.025000 0.725000 1.755000 0.895000 ;
        RECT 1.045000 1.630000 1.235000 2.435000 ;
        RECT 1.475000 0.895000 1.755000 1.460000 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.800000 0.875000 2.465000 ;
      LAYER mcon ;
        RECT 0.600000 2.125000 0.770000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.405000 1.800000 1.735000 2.465000 ;
      LAYER mcon ;
        RECT 1.500000 2.125000 1.670000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 1.770000 2.340000 ;
        RECT 0.540000 2.080000 0.830000 2.140000 ;
        RECT 1.440000 2.080000 1.730000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.560000  0.085000 0.855000 0.610000 ;
      RECT 1.420000  0.085000 1.750000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_2
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  4.608000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.345000 0.895000  2.155000 1.275000 ;
        RECT 8.930000 0.895000 10.710000 1.275000 ;
      LAYER mcon ;
        RECT 1.525000 1.105000 1.695000 1.275000 ;
        RECT 1.985000 1.105000 2.155000 1.275000 ;
        RECT 9.345000 1.105000 9.515000 1.275000 ;
        RECT 9.805000 1.105000 9.975000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465000 1.075000  2.215000 1.120000 ;
        RECT 1.465000 1.120000 10.035000 1.260000 ;
        RECT 1.465000 1.260000  2.215000 1.305000 ;
        RECT 9.285000 1.075000 10.035000 1.120000 ;
        RECT 9.285000 1.260000 10.035000 1.305000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.520900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.615000 1.455000 10.480000 1.665000 ;
        RECT  0.615000 1.665000  0.785000 2.465000 ;
        RECT  1.475000 1.665000  1.645000 2.465000 ;
        RECT  2.325000 0.280000  2.550000 1.415000 ;
        RECT  2.325000 1.415000  8.755000 1.455000 ;
        RECT  2.335000 1.665000  2.505000 2.465000 ;
        RECT  3.155000 0.280000  3.410000 1.415000 ;
        RECT  3.195000 1.665000  3.365000 2.465000 ;
        RECT  4.015000 0.280000  4.255000 1.415000 ;
        RECT  4.055000 1.665000  4.225000 2.465000 ;
        RECT  4.905000 0.280000  5.255000 1.415000 ;
        RECT  5.080000 1.665000  5.250000 2.465000 ;
        RECT  5.925000 0.280000  6.175000 1.415000 ;
        RECT  5.965000 1.665000  6.135000 2.465000 ;
        RECT  6.785000 0.280000  7.035000 1.415000 ;
        RECT  6.825000 1.665000  6.995000 2.465000 ;
        RECT  7.645000 0.280000  7.895000 1.415000 ;
        RECT  7.685000 1.665000  7.855000 2.465000 ;
        RECT  8.505000 0.280000  8.755000 1.415000 ;
        RECT  8.545000 1.665000  8.715000 2.465000 ;
        RECT  9.405000 1.665000  9.575000 2.465000 ;
        RECT 10.265000 1.665000 10.435000 2.465000 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.110000 1.495000  0.440000 2.465000 ;
        RECT 10.610000 1.835000 10.940000 2.465000 ;
      LAYER mcon ;
        RECT  0.130000 2.125000  0.300000 2.295000 ;
        RECT 10.720000 2.125000 10.890000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.965000 1.835000 1.295000 2.465000 ;
      LAYER mcon ;
        RECT 0.990000 2.125000 1.160000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.825000 1.835000 2.155000 2.465000 ;
      LAYER mcon ;
        RECT 1.890000 2.125000 2.060000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.685000 1.835000 3.015000 2.465000 ;
      LAYER mcon ;
        RECT 2.770000 2.125000 2.940000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.545000 1.835000 3.875000 2.465000 ;
      LAYER mcon ;
        RECT 3.690000 2.125000 3.860000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.425000 1.835000 4.755000 2.465000 ;
      LAYER mcon ;
        RECT 4.550000 2.125000 4.720000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.450000 1.835000 5.780000 2.465000 ;
      LAYER mcon ;
        RECT 5.450000 2.125000 5.620000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.315000 1.835000 6.645000 2.465000 ;
      LAYER mcon ;
        RECT 6.370000 2.125000 6.540000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.175000 1.835000 7.505000 2.465000 ;
      LAYER mcon ;
        RECT 7.230000 2.125000 7.400000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.035000 1.835000 8.365000 2.465000 ;
      LAYER mcon ;
        RECT 8.130000 2.125000 8.300000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.895000 1.835000 9.225000 2.465000 ;
      LAYER mcon ;
        RECT 8.960000 2.125000 9.130000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755000 1.835000 10.085000 2.465000 ;
      LAYER mcon ;
        RECT 9.820000 2.125000 9.990000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT  0.070000 2.080000  0.360000 2.140000 ;
        RECT  0.070000 2.140000 10.970000 2.340000 ;
        RECT  0.930000 2.080000  1.220000 2.140000 ;
        RECT  1.830000 2.080000  2.120000 2.140000 ;
        RECT  2.710000 2.080000  3.000000 2.140000 ;
        RECT  3.630000 2.080000  3.920000 2.140000 ;
        RECT  4.490000 2.080000  4.780000 2.140000 ;
        RECT  5.390000 2.080000  5.680000 2.140000 ;
        RECT  6.310000 2.080000  6.600000 2.140000 ;
        RECT  7.170000 2.080000  7.460000 2.140000 ;
        RECT  8.070000 2.080000  8.360000 2.140000 ;
        RECT  8.900000 2.080000  9.190000 2.140000 ;
        RECT  9.760000 2.080000 10.050000 2.140000 ;
        RECT 10.660000 2.080000 10.950000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 11.040000 0.085000 ;
      RECT 0.000000  2.635000 11.040000 2.805000 ;
      RECT 1.855000  0.085000  2.125000 0.610000 ;
      RECT 2.720000  0.085000  2.985000 0.610000 ;
      RECT 3.580000  0.085000  3.845000 0.610000 ;
      RECT 4.465000  0.085000  4.730000 0.610000 ;
      RECT 5.490000  0.085000  5.755000 0.610000 ;
      RECT 6.350000  0.085000  6.575000 0.610000 ;
      RECT 7.210000  0.085000  7.475000 0.610000 ;
      RECT 8.070000  0.085000  8.335000 0.610000 ;
      RECT 8.930000  0.085000  9.195000 0.610000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_16
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.304000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.035000 4.865000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.090400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.695000 5.440000 0.865000 ;
        RECT 0.115000 0.865000 0.285000 1.460000 ;
        RECT 0.115000 1.460000 5.440000 1.630000 ;
        RECT 0.595000 1.630000 0.765000 2.435000 ;
        RECT 1.440000 1.630000 1.610000 2.435000 ;
        RECT 1.535000 0.280000 1.725000 0.695000 ;
        RECT 2.280000 1.630000 2.450000 2.435000 ;
        RECT 2.395000 0.280000 2.585000 0.695000 ;
        RECT 3.120000 1.630000 3.290000 2.435000 ;
        RECT 3.255000 0.280000 3.445000 0.695000 ;
        RECT 3.960000 1.630000 4.130000 2.435000 ;
        RECT 4.115000 0.280000 4.305000 0.695000 ;
        RECT 4.800000 1.630000 4.970000 2.435000 ;
        RECT 5.170000 0.865000 5.440000 1.460000 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.800000 0.425000 2.465000 ;
        RECT 5.140000 1.800000 5.470000 2.465000 ;
      LAYER mcon ;
        RECT 0.130000 2.125000 0.300000 2.295000 ;
        RECT 5.255000 2.125000 5.425000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.940000 1.800000 1.270000 2.465000 ;
      LAYER mcon ;
        RECT 0.990000 2.125000 1.160000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.780000 1.800000 2.110000 2.465000 ;
      LAYER mcon ;
        RECT 1.890000 2.125000 2.060000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.620000 1.800000 2.950000 2.465000 ;
      LAYER mcon ;
        RECT 2.770000 2.125000 2.940000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.460000 1.800000 3.790000 2.465000 ;
      LAYER mcon ;
        RECT 3.495000 2.125000 3.665000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.300000 1.800000 4.630000 2.465000 ;
      LAYER mcon ;
        RECT 4.355000 2.125000 4.525000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.080000 0.360000 2.140000 ;
        RECT 0.070000 2.140000 5.910000 2.340000 ;
        RECT 0.930000 2.080000 1.220000 2.140000 ;
        RECT 1.830000 2.080000 2.120000 2.140000 ;
        RECT 2.710000 2.080000 3.000000 2.140000 ;
        RECT 3.435000 2.080000 3.725000 2.140000 ;
        RECT 4.295000 2.080000 4.585000 2.140000 ;
        RECT 5.195000 2.080000 5.485000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 1.035000  0.085000 1.365000 0.525000 ;
      RECT 1.895000  0.085000 2.225000 0.525000 ;
      RECT 2.755000  0.085000 3.085000 0.525000 ;
      RECT 3.615000  0.085000 3.945000 0.525000 ;
      RECT 4.475000  0.085000 4.805000 0.525000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_8
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.375000 0.325000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.336000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 0.255000 0.840000 0.760000 ;
        RECT 0.590000 0.760000 1.295000 0.945000 ;
        RECT 0.595000 0.945000 1.295000 1.290000 ;
        RECT 0.595000 1.290000 0.765000 2.465000 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.665000 0.425000 2.465000 ;
      LAYER mcon ;
        RECT 0.155000 2.125000 0.325000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.935000 1.665000 1.295000 2.465000 ;
      LAYER mcon ;
        RECT 1.055000 2.125000 1.225000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 1.310000 2.340000 ;
        RECT 0.095000 2.080000 0.385000 2.140000 ;
        RECT 0.995000 2.080000 1.285000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 1.010000  0.085000 1.295000 0.590000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_1
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.152000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.065000 2.660000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.075200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.725000 3.135000 0.895000 ;
        RECT 0.105000 0.895000 0.275000 1.460000 ;
        RECT 0.105000 1.460000 3.135000 1.630000 ;
        RECT 0.645000 1.630000 0.815000 2.435000 ;
        RECT 1.030000 0.280000 1.290000 0.725000 ;
        RECT 1.505000 1.630000 1.675000 2.435000 ;
        RECT 1.890000 0.280000 2.145000 0.725000 ;
        RECT 2.365000 1.630000 2.535000 2.435000 ;
        RECT 2.835000 0.895000 3.135000 1.460000 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.135000 1.800000 0.465000 2.465000 ;
      LAYER mcon ;
        RECT 0.195000 2.125000 0.365000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.995000 1.800000 1.325000 2.465000 ;
      LAYER mcon ;
        RECT 1.055000 2.125000 1.225000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.855000 1.800000 2.185000 2.465000 ;
      LAYER mcon ;
        RECT 1.955000 2.125000 2.125000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.715000 1.800000 3.045000 2.465000 ;
      LAYER mcon ;
        RECT 2.835000 2.125000 3.005000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 3.150000 2.340000 ;
        RECT 0.135000 2.080000 0.425000 2.140000 ;
        RECT 0.995000 2.080000 1.285000 2.140000 ;
        RECT 1.895000 2.080000 2.185000 2.140000 ;
        RECT 2.775000 2.080000 3.065000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.565000  0.085000 0.860000 0.555000 ;
      RECT 1.460000  0.085000 1.720000 0.555000 ;
      RECT 2.315000  0.085000 2.615000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_4
MACRO sky130_fd_sc_hd__and2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.445000 1.615000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 1.645000 2.175000 1.955000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.350000 1.580000 2.655000 2.365000 ;
        RECT 2.415000 0.255000 2.655000 0.775000 ;
        RECT 2.480000 0.775000 2.655000 1.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.590000 ;
      RECT 0.175000  1.785000 0.850000 2.015000 ;
      RECT 0.175000  2.015000 0.345000 2.445000 ;
      RECT 0.515000  2.185000 0.845000 2.635000 ;
      RECT 0.595000  0.280000 0.835000 0.655000 ;
      RECT 0.615000  0.655000 0.835000 0.805000 ;
      RECT 0.615000  0.805000 1.150000 1.135000 ;
      RECT 0.615000  1.135000 0.850000 1.785000 ;
      RECT 1.020000  1.305000 2.305000 1.325000 ;
      RECT 1.020000  1.325000 1.880000 1.475000 ;
      RECT 1.020000  1.475000 1.305000 2.420000 ;
      RECT 1.115000  0.270000 1.285000 0.415000 ;
      RECT 1.115000  0.415000 1.490000 0.610000 ;
      RECT 1.320000  0.610000 1.490000 0.945000 ;
      RECT 1.320000  0.945000 2.305000 1.305000 ;
      RECT 1.485000  2.165000 2.170000 2.635000 ;
      RECT 1.850000  0.085000 2.245000 0.580000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__and2b_1
MACRO sky130_fd_sc_hd__and2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.900000 0.625000 3.155000 0.995000 ;
        RECT 2.900000 0.995000 3.205000 1.325000 ;
        RECT 2.900000 1.325000 3.155000 1.745000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 0.995000 0.975000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.934000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.535000 2.730000 1.745000 ;
        RECT 1.525000 0.495000 1.715000 0.615000 ;
        RECT 1.525000 0.615000 2.730000 0.825000 ;
        RECT 2.440000 0.825000 2.730000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.615000 ;
      RECT 0.090000  0.615000 1.355000 0.805000 ;
      RECT 0.090000  2.255000 0.425000 2.635000 ;
      RECT 0.165000  0.995000 0.425000 1.325000 ;
      RECT 0.165000  1.325000 0.335000 1.915000 ;
      RECT 0.165000  1.915000 3.505000 2.085000 ;
      RECT 0.515000  1.500000 1.315000 1.745000 ;
      RECT 0.955000  0.085000 1.285000 0.445000 ;
      RECT 0.990000  2.275000 1.320000 2.635000 ;
      RECT 1.110000  1.435000 1.320000 1.485000 ;
      RECT 1.110000  1.485000 1.315000 1.500000 ;
      RECT 1.145000  0.805000 1.355000 0.995000 ;
      RECT 1.145000  0.995000 2.260000 1.355000 ;
      RECT 1.145000  1.355000 1.320000 1.435000 ;
      RECT 1.885000  0.085000 2.215000 0.445000 ;
      RECT 1.905000  2.275000 2.235000 2.635000 ;
      RECT 2.745000  0.085000 3.075000 0.445000 ;
      RECT 2.745000  2.275000 3.075000 2.635000 ;
      RECT 3.330000  0.495000 3.500000 0.675000 ;
      RECT 3.330000  0.675000 3.545000 0.845000 ;
      RECT 3.335000  1.530000 3.545000 1.700000 ;
      RECT 3.335000  1.700000 3.505000 1.915000 ;
      RECT 3.375000  0.845000 3.545000 1.530000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__and2b_4
MACRO sky130_fd_sc_hd__and2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.765000 0.450000 1.615000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.645000 2.200000 1.955000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 1.580000 2.680000 2.365000 ;
        RECT 2.445000 0.255000 2.680000 0.775000 ;
        RECT 2.505000 0.775000 2.680000 1.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.590000 ;
      RECT 0.175000  1.785000 0.855000 2.015000 ;
      RECT 0.175000  2.015000 0.345000 2.445000 ;
      RECT 0.515000  2.185000 0.845000 2.635000 ;
      RECT 0.595000  0.280000 0.835000 0.655000 ;
      RECT 0.620000  0.655000 0.835000 0.805000 ;
      RECT 0.620000  0.805000 1.175000 1.135000 ;
      RECT 0.620000  1.135000 0.855000 1.785000 ;
      RECT 1.045000  1.305000 2.335000 1.325000 ;
      RECT 1.045000  1.325000 1.905000 1.475000 ;
      RECT 1.045000  1.475000 1.330000 2.420000 ;
      RECT 1.115000  0.270000 1.285000 0.415000 ;
      RECT 1.115000  0.415000 1.515000 0.610000 ;
      RECT 1.345000  0.610000 1.515000 0.945000 ;
      RECT 1.345000  0.945000 2.335000 1.305000 ;
      RECT 1.510000  2.165000 2.195000 2.635000 ;
      RECT 1.875000  0.085000 2.275000 0.580000 ;
      RECT 2.865000  0.085000 3.135000 0.720000 ;
      RECT 2.865000  1.680000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__and2b_2
MACRO sky130_fd_sc_hd__dlymetal6s6s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s6s_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.575000 1.700000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.080000 0.255000 4.515000 0.825000 ;
        RECT 4.080000 1.495000 4.515000 2.465000 ;
        RECT 4.155000 0.825000 4.515000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125000 -0.085000 0.295000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.255000 0.525000 0.655000 ;
      RECT 0.085000  0.655000 1.080000 0.825000 ;
      RECT 0.085000  1.870000 1.080000 2.040000 ;
      RECT 0.085000  2.040000 0.525000 2.465000 ;
      RECT 0.695000  0.085000 1.080000 0.485000 ;
      RECT 0.695000  2.210000 1.080000 2.635000 ;
      RECT 0.745000  0.825000 1.080000 0.995000 ;
      RECT 0.745000  0.995000 1.155000 1.325000 ;
      RECT 0.745000  1.325000 1.080000 1.870000 ;
      RECT 1.250000  0.255000 1.520000 0.825000 ;
      RECT 1.250000  1.495000 1.975000 1.675000 ;
      RECT 1.250000  1.675000 1.520000 2.465000 ;
      RECT 1.325000  0.825000 1.520000 0.995000 ;
      RECT 1.325000  0.995000 1.975000 1.495000 ;
      RECT 1.690000  0.255000 1.940000 0.655000 ;
      RECT 1.690000  0.655000 2.495000 0.825000 ;
      RECT 1.690000  1.845000 2.495000 2.040000 ;
      RECT 1.690000  2.040000 1.940000 2.465000 ;
      RECT 2.110000  0.085000 2.495000 0.485000 ;
      RECT 2.110000  2.210000 2.495000 2.635000 ;
      RECT 2.145000  0.825000 2.495000 0.995000 ;
      RECT 2.145000  0.995000 2.570000 1.325000 ;
      RECT 2.145000  1.325000 2.495000 1.845000 ;
      RECT 2.665000  0.255000 2.915000 0.825000 ;
      RECT 2.665000  1.495000 3.390000 1.675000 ;
      RECT 2.665000  1.675000 2.915000 2.465000 ;
      RECT 2.740000  0.825000 2.915000 0.995000 ;
      RECT 2.740000  0.995000 3.390000 1.495000 ;
      RECT 3.085000  0.255000 3.355000 0.655000 ;
      RECT 3.085000  0.655000 3.910000 0.825000 ;
      RECT 3.085000  1.845000 3.910000 2.040000 ;
      RECT 3.085000  2.040000 3.355000 2.465000 ;
      RECT 3.525000  0.085000 3.910000 0.485000 ;
      RECT 3.525000  2.210000 3.910000 2.635000 ;
      RECT 3.560000  0.825000 3.910000 0.995000 ;
      RECT 3.560000  0.995000 3.985000 1.325000 ;
      RECT 3.560000  1.325000 3.910000 1.845000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__dlymetal6s6s_1
MACRO sky130_fd_sc_hd__lpflow_inputiso1n_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso1n_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 2.085000 1.735000 2.415000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.325000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 0.415000 2.675000 0.760000 ;
        RECT 2.405000 1.495000 2.675000 2.465000 ;
        RECT 2.505000 0.760000 2.675000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.110000  0.265000 0.420000 0.735000 ;
      RECT 0.110000  0.735000 0.845000 0.905000 ;
      RECT 0.590000  0.085000 1.325000 0.565000 ;
      RECT 0.595000  0.905000 0.845000 0.995000 ;
      RECT 0.595000  0.995000 1.335000 1.325000 ;
      RECT 0.595000  1.325000 0.765000 1.885000 ;
      RECT 0.990000  1.495000 2.235000 1.665000 ;
      RECT 0.990000  1.665000 1.410000 1.915000 ;
      RECT 1.495000  0.305000 1.665000 0.655000 ;
      RECT 1.495000  0.655000 2.235000 0.825000 ;
      RECT 1.835000  0.085000 2.215000 0.485000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
      RECT 2.065000  0.825000 2.235000 0.995000 ;
      RECT 2.065000  0.995000 2.295000 1.325000 ;
      RECT 2.065000  1.325000 2.235000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso1n_1
MACRO sky130_fd_sc_hd__dlxbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 0.955000 1.810000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.215000 0.415000 5.465000 0.660000 ;
        RECT 5.215000 0.660000 5.500000 0.825000 ;
        RECT 5.215000 1.495000 5.500000 1.710000 ;
        RECT 5.215000 1.710000 5.465000 2.455000 ;
        RECT 5.330000 0.825000 5.500000 0.995000 ;
        RECT 5.330000 0.995000 5.905000 1.325000 ;
        RECT 5.330000 1.325000 5.500000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.050000 0.255000 7.305000 0.825000 ;
        RECT 7.050000 1.445000 7.305000 2.465000 ;
        RECT 7.095000 0.825000 7.305000 1.055000 ;
        RECT 7.095000 1.055000 7.735000 1.325000 ;
        RECT 7.095000 1.325000 7.305000 1.445000 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.475000  1.495000 2.160000 1.665000 ;
      RECT 1.475000  1.665000 1.805000 2.415000 ;
      RECT 1.555000  0.345000 1.725000 0.615000 ;
      RECT 1.555000  0.615000 2.160000 0.765000 ;
      RECT 1.555000  0.765000 2.360000 0.785000 ;
      RECT 1.895000  0.085000 2.225000 0.445000 ;
      RECT 1.975000  1.835000 2.290000 2.635000 ;
      RECT 1.990000  0.785000 2.360000 1.095000 ;
      RECT 1.990000  1.095000 2.160000 1.495000 ;
      RECT 2.490000  1.355000 2.775000 2.005000 ;
      RECT 2.735000  0.705000 3.115000 1.035000 ;
      RECT 2.860000  0.365000 3.520000 0.535000 ;
      RECT 2.920000  2.255000 3.670000 2.425000 ;
      RECT 2.945000  1.035000 3.115000 1.415000 ;
      RECT 2.945000  1.415000 3.285000 1.995000 ;
      RECT 3.350000  0.535000 3.520000 0.995000 ;
      RECT 3.350000  0.995000 4.220000 1.165000 ;
      RECT 3.500000  1.165000 4.220000 1.325000 ;
      RECT 3.500000  1.325000 3.670000 2.255000 ;
      RECT 3.760000  0.085000 4.090000 0.825000 ;
      RECT 3.840000  2.135000 4.140000 2.635000 ;
      RECT 3.860000  1.535000 4.580000 1.865000 ;
      RECT 4.360000  0.415000 4.580000 0.825000 ;
      RECT 4.360000  1.865000 4.580000 2.435000 ;
      RECT 4.410000  0.825000 4.580000 0.995000 ;
      RECT 4.410000  0.995000 5.160000 1.325000 ;
      RECT 4.410000  1.325000 4.580000 1.535000 ;
      RECT 4.760000  0.085000 5.045000 0.825000 ;
      RECT 4.760000  1.495000 5.045000 2.635000 ;
      RECT 5.635000  0.085000 5.905000 0.545000 ;
      RECT 5.635000  1.835000 5.905000 2.635000 ;
      RECT 6.075000  0.255000 6.405000 0.995000 ;
      RECT 6.075000  0.995000 6.925000 1.325000 ;
      RECT 6.075000  1.325000 6.405000 2.465000 ;
      RECT 6.585000  0.085000 6.880000 0.545000 ;
      RECT 6.585000  1.835000 6.880000 2.635000 ;
      RECT 7.475000  0.085000 7.735000 0.885000 ;
      RECT 7.475000  1.495000 7.735000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.490000  1.785000 2.660000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.950000  1.445000 3.120000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.180000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.720000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.430000 1.755000 2.720000 1.800000 ;
      RECT 2.430000 1.940000 2.720000 1.985000 ;
      RECT 2.890000 1.415000 3.180000 1.460000 ;
      RECT 2.890000 1.600000 3.180000 1.645000 ;
  END
END sky130_fd_sc_hd__dlxbn_2
MACRO sky130_fd_sc_hd__dlxbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 0.955000 1.785000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.140000 0.415000 5.480000 0.745000 ;
        RECT 5.140000 1.670000 5.480000 2.465000 ;
        RECT 5.310000 0.745000 5.480000 1.670000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.555000 0.255000 6.815000 0.825000 ;
        RECT 6.555000 1.505000 6.815000 2.465000 ;
        RECT 6.625000 0.825000 6.815000 1.505000 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.480000  1.495000 2.165000 1.665000 ;
      RECT 1.480000  1.665000 1.810000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.165000 0.785000 ;
      RECT 1.875000  0.085000 2.230000 0.445000 ;
      RECT 1.980000  1.835000 2.295000 2.635000 ;
      RECT 1.995000  0.785000 2.165000 0.905000 ;
      RECT 1.995000  0.905000 2.365000 1.235000 ;
      RECT 1.995000  1.235000 2.165000 1.495000 ;
      RECT 2.495000  1.355000 2.780000 2.005000 ;
      RECT 2.565000  0.705000 3.120000 1.035000 ;
      RECT 2.790000  0.365000 3.525000 0.535000 ;
      RECT 2.920000  2.105000 3.620000 2.115000 ;
      RECT 2.920000  2.115000 3.615000 2.130000 ;
      RECT 2.920000  2.130000 3.610000 2.275000 ;
      RECT 2.950000  1.035000 3.120000 1.415000 ;
      RECT 2.950000  1.415000 3.290000 1.910000 ;
      RECT 3.355000  0.535000 3.525000 0.995000 ;
      RECT 3.355000  0.995000 4.225000 1.165000 ;
      RECT 3.360000  2.075000 3.630000 2.090000 ;
      RECT 3.360000  2.090000 3.625000 2.105000 ;
      RECT 3.375000  2.060000 3.630000 2.075000 ;
      RECT 3.420000  2.030000 3.630000 2.060000 ;
      RECT 3.430000  2.015000 3.630000 2.030000 ;
      RECT 3.460000  1.165000 4.225000 1.325000 ;
      RECT 3.460000  1.325000 3.630000 2.015000 ;
      RECT 3.765000  0.085000 4.095000 0.610000 ;
      RECT 3.780000  2.175000 3.950000 2.635000 ;
      RECT 3.800000  1.535000 4.580000 1.620000 ;
      RECT 3.800000  1.620000 4.550000 1.865000 ;
      RECT 4.300000  0.415000 4.470000 0.660000 ;
      RECT 4.300000  0.660000 4.580000 0.840000 ;
      RECT 4.300000  1.865000 4.550000 2.435000 ;
      RECT 4.395000  0.840000 4.580000 0.995000 ;
      RECT 4.395000  0.995000 5.140000 1.325000 ;
      RECT 4.395000  1.325000 4.580000 1.535000 ;
      RECT 4.640000  0.085000 4.970000 0.495000 ;
      RECT 4.720000  1.830000 4.970000 2.635000 ;
      RECT 5.660000  0.255000 5.910000 0.995000 ;
      RECT 5.660000  0.995000 6.455000 1.325000 ;
      RECT 5.660000  1.325000 5.910000 2.465000 ;
      RECT 6.090000  0.085000 6.385000 0.545000 ;
      RECT 6.090000  1.835000 6.385000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.495000  1.785000 2.665000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.955000  1.445000 3.125000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.185000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.725000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.435000 1.755000 2.725000 1.800000 ;
      RECT 2.435000 1.940000 2.725000 1.985000 ;
      RECT 2.895000 1.415000 3.185000 1.460000 ;
      RECT 2.895000 1.600000 3.185000 1.645000 ;
  END
END sky130_fd_sc_hd__dlxbn_1
MACRO sky130_fd_sc_hd__dfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 1.065000 1.720000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.985000 0.305000 7.320000 0.730000 ;
        RECT 6.985000 0.730000 8.655000 0.900000 ;
        RECT 6.985000 1.465000 8.655000 1.635000 ;
        RECT 6.985000 1.635000 7.320000 2.395000 ;
        RECT 7.840000 0.305000 8.175000 0.730000 ;
        RECT 7.840000 1.635000 8.170000 2.395000 ;
        RECT 8.410000 0.900000 8.655000 1.465000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.240000 2.465000 ;
      RECT 1.440000  2.175000 1.705000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.890000  0.365000 2.220000 0.535000 ;
      RECT 1.890000  0.535000 2.060000 2.065000 ;
      RECT 1.890000  2.065000 2.125000 2.440000 ;
      RECT 2.230000  0.705000 2.810000 1.035000 ;
      RECT 2.230000  1.035000 2.470000 1.905000 ;
      RECT 2.370000  2.190000 3.440000 2.360000 ;
      RECT 2.400000  0.365000 3.150000 0.535000 ;
      RECT 2.660000  1.655000 3.100000 2.010000 ;
      RECT 2.980000  0.535000 3.150000 1.315000 ;
      RECT 2.980000  1.315000 3.780000 1.485000 ;
      RECT 3.270000  1.485000 3.780000 1.575000 ;
      RECT 3.270000  1.575000 3.440000 2.190000 ;
      RECT 3.320000  0.765000 4.120000 1.065000 ;
      RECT 3.320000  1.065000 3.490000 1.095000 ;
      RECT 3.400000  0.085000 3.770000 0.585000 ;
      RECT 3.610000  1.245000 3.780000 1.315000 ;
      RECT 3.610000  1.835000 3.780000 2.635000 ;
      RECT 3.950000  0.365000 4.410000 0.535000 ;
      RECT 3.950000  0.535000 4.120000 0.765000 ;
      RECT 3.950000  1.065000 4.120000 2.135000 ;
      RECT 3.950000  2.135000 4.200000 2.465000 ;
      RECT 4.290000  0.705000 4.840000 1.035000 ;
      RECT 4.290000  1.245000 4.480000 1.965000 ;
      RECT 4.425000  2.165000 5.310000 2.335000 ;
      RECT 4.640000  0.365000 5.310000 0.535000 ;
      RECT 4.650000  1.035000 4.840000 1.575000 ;
      RECT 4.650000  1.575000 4.970000 1.905000 ;
      RECT 5.140000  0.535000 5.310000 1.075000 ;
      RECT 5.140000  1.075000 6.230000 1.245000 ;
      RECT 5.140000  1.245000 5.310000 2.165000 ;
      RECT 5.480000  1.500000 6.590000 1.670000 ;
      RECT 5.480000  1.670000 6.340000 1.830000 ;
      RECT 5.490000  2.135000 5.705000 2.635000 ;
      RECT 5.625000  0.085000 5.795000 0.615000 ;
      RECT 6.090000  0.295000 6.450000 0.735000 ;
      RECT 6.090000  0.735000 6.590000 0.905000 ;
      RECT 6.170000  1.830000 6.340000 2.455000 ;
      RECT 6.420000  0.905000 6.590000 1.075000 ;
      RECT 6.420000  1.075000 8.240000 1.245000 ;
      RECT 6.420000  1.245000 6.590000 1.500000 ;
      RECT 6.625000  0.085000 6.795000 0.565000 ;
      RECT 6.625000  1.855000 6.805000 2.635000 ;
      RECT 7.495000  0.085000 7.665000 0.560000 ;
      RECT 7.500000  1.805000 7.670000 2.635000 ;
      RECT 8.340000  1.805000 8.510000 2.635000 ;
      RECT 8.345000  0.085000 8.515000 0.560000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.785000 0.780000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  0.765000 1.240000 0.935000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  0.765000 2.640000 0.935000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.785000 3.100000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.310000  0.765000 4.480000 0.935000 ;
      RECT 4.310000  1.785000 4.480000 1.955000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.755000 0.840000 1.800000 ;
      RECT 0.550000 1.800000 4.540000 1.940000 ;
      RECT 0.550000 1.940000 0.840000 1.985000 ;
      RECT 1.010000 0.735000 1.300000 0.780000 ;
      RECT 1.010000 0.780000 4.540000 0.920000 ;
      RECT 1.010000 0.920000 1.300000 0.965000 ;
      RECT 2.410000 0.735000 2.700000 0.780000 ;
      RECT 2.410000 0.920000 2.700000 0.965000 ;
      RECT 2.870000 1.755000 3.160000 1.800000 ;
      RECT 2.870000 1.940000 3.160000 1.985000 ;
      RECT 4.250000 0.735000 4.540000 0.780000 ;
      RECT 4.250000 0.920000 4.540000 0.965000 ;
      RECT 4.250000 1.755000 4.540000 1.800000 ;
      RECT 4.250000 1.940000 4.540000 1.985000 ;
  END
END sky130_fd_sc_hd__dfxtp_4
MACRO sky130_fd_sc_hd__dfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.370000 0.715000 1.650000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.885000 1.495000 7.275000 1.575000 ;
        RECT 6.885000 1.575000 7.215000 2.420000 ;
        RECT 6.895000 0.305000 7.225000 0.740000 ;
        RECT 6.895000 0.740000 7.275000 0.825000 ;
        RECT 7.050000 0.825000 7.275000 0.865000 ;
        RECT 7.060000 1.445000 7.275000 1.495000 ;
        RECT 7.105000 0.865000 7.275000 1.445000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.200000 2.465000 ;
      RECT 1.440000  2.175000 1.705000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.820000  0.675000 2.045000 0.805000 ;
      RECT 1.820000  0.805000 1.990000 1.910000 ;
      RECT 1.820000  1.910000 2.125000 2.040000 ;
      RECT 1.875000  0.365000 2.210000 0.535000 ;
      RECT 1.875000  0.535000 2.045000 0.675000 ;
      RECT 1.875000  2.040000 2.125000 2.465000 ;
      RECT 2.160000  1.125000 2.400000 1.720000 ;
      RECT 2.215000  0.735000 2.740000 0.955000 ;
      RECT 2.335000  2.190000 3.440000 2.360000 ;
      RECT 2.405000  0.365000 3.080000 0.535000 ;
      RECT 2.570000  0.955000 2.740000 1.655000 ;
      RECT 2.570000  1.655000 3.100000 2.020000 ;
      RECT 2.910000  0.535000 3.080000 1.315000 ;
      RECT 2.910000  1.315000 3.780000 1.485000 ;
      RECT 3.270000  1.485000 3.780000 1.575000 ;
      RECT 3.270000  1.575000 3.440000 2.190000 ;
      RECT 3.290000  0.765000 4.120000 1.065000 ;
      RECT 3.290000  1.065000 3.490000 1.095000 ;
      RECT 3.400000  0.085000 3.770000 0.585000 ;
      RECT 3.610000  1.245000 3.780000 1.315000 ;
      RECT 3.610000  1.835000 3.780000 2.635000 ;
      RECT 3.950000  0.365000 4.355000 0.535000 ;
      RECT 3.950000  0.535000 4.120000 0.765000 ;
      RECT 3.950000  1.065000 4.120000 2.135000 ;
      RECT 3.950000  2.135000 4.200000 2.465000 ;
      RECT 4.290000  1.245000 4.480000 1.965000 ;
      RECT 4.425000  2.165000 5.310000 2.335000 ;
      RECT 4.505000  0.705000 4.970000 1.035000 ;
      RECT 4.525000  0.365000 5.310000 0.535000 ;
      RECT 4.650000  1.035000 4.970000 1.995000 ;
      RECT 5.140000  0.535000 5.310000 0.995000 ;
      RECT 5.140000  0.995000 6.015000 1.325000 ;
      RECT 5.140000  1.325000 5.310000 2.165000 ;
      RECT 5.480000  1.530000 6.375000 1.905000 ;
      RECT 5.490000  2.135000 5.805000 2.635000 ;
      RECT 5.585000  0.085000 5.795000 0.615000 ;
      RECT 6.035000  1.905000 6.375000 2.465000 ;
      RECT 6.055000  0.300000 6.385000 0.825000 ;
      RECT 6.185000  0.825000 6.385000 0.995000 ;
      RECT 6.185000  0.995000 6.935000 1.325000 ;
      RECT 6.185000  1.325000 6.375000 1.530000 ;
      RECT 6.545000  1.625000 6.715000 2.635000 ;
      RECT 6.555000  0.085000 6.725000 0.695000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.630000  1.785000 0.800000 1.955000 ;
      RECT 1.025000  1.445000 1.195000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.215000  1.445000 2.385000 1.615000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.730000  1.785000 2.900000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.300000  1.785000 4.470000 1.955000 ;
      RECT 4.735000  1.445000 4.905000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 0.570000 1.755000 0.860000 1.800000 ;
      RECT 0.570000 1.800000 4.530000 1.940000 ;
      RECT 0.570000 1.940000 0.860000 1.985000 ;
      RECT 0.965000 1.415000 1.255000 1.460000 ;
      RECT 0.965000 1.460000 4.965000 1.600000 ;
      RECT 0.965000 1.600000 1.255000 1.645000 ;
      RECT 2.155000 1.415000 2.445000 1.460000 ;
      RECT 2.155000 1.600000 2.445000 1.645000 ;
      RECT 2.670000 1.755000 2.960000 1.800000 ;
      RECT 2.670000 1.940000 2.960000 1.985000 ;
      RECT 4.240000 1.755000 4.530000 1.800000 ;
      RECT 4.240000 1.940000 4.530000 1.985000 ;
      RECT 4.675000 1.415000 4.965000 1.460000 ;
      RECT 4.675000 1.600000 4.965000 1.645000 ;
  END
END sky130_fd_sc_hd__dfxtp_1
MACRO sky130_fd_sc_hd__dfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.370000 0.715000 1.650000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.885000 1.495000 7.275000 1.575000 ;
        RECT 6.885000 1.575000 7.215000 2.420000 ;
        RECT 6.895000 0.305000 7.225000 0.740000 ;
        RECT 6.895000 0.740000 7.275000 0.825000 ;
        RECT 7.050000 0.825000 7.275000 0.865000 ;
        RECT 7.060000 1.445000 7.275000 1.495000 ;
        RECT 7.105000 0.865000 7.275000 1.445000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.200000 2.465000 ;
      RECT 1.440000  2.175000 1.705000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.820000  0.675000 2.045000 0.805000 ;
      RECT 1.820000  0.805000 1.990000 1.910000 ;
      RECT 1.820000  1.910000 2.125000 2.040000 ;
      RECT 1.875000  0.365000 2.210000 0.535000 ;
      RECT 1.875000  0.535000 2.045000 0.675000 ;
      RECT 1.875000  2.040000 2.125000 2.465000 ;
      RECT 2.160000  1.125000 2.400000 1.720000 ;
      RECT 2.215000  0.735000 2.740000 0.955000 ;
      RECT 2.335000  2.190000 3.440000 2.360000 ;
      RECT 2.405000  0.365000 3.080000 0.535000 ;
      RECT 2.570000  0.955000 2.740000 1.655000 ;
      RECT 2.570000  1.655000 3.100000 2.020000 ;
      RECT 2.910000  0.535000 3.080000 1.315000 ;
      RECT 2.910000  1.315000 3.780000 1.485000 ;
      RECT 3.270000  1.485000 3.780000 1.575000 ;
      RECT 3.270000  1.575000 3.440000 2.190000 ;
      RECT 3.290000  0.765000 4.120000 1.065000 ;
      RECT 3.290000  1.065000 3.490000 1.095000 ;
      RECT 3.400000  0.085000 3.770000 0.585000 ;
      RECT 3.610000  1.245000 3.780000 1.315000 ;
      RECT 3.610000  1.835000 3.780000 2.635000 ;
      RECT 3.950000  0.365000 4.355000 0.535000 ;
      RECT 3.950000  0.535000 4.120000 0.765000 ;
      RECT 3.950000  1.065000 4.120000 2.135000 ;
      RECT 3.950000  2.135000 4.200000 2.465000 ;
      RECT 4.290000  1.245000 4.480000 1.965000 ;
      RECT 4.425000  2.165000 5.310000 2.335000 ;
      RECT 4.505000  0.705000 4.970000 1.035000 ;
      RECT 4.525000  0.365000 5.310000 0.535000 ;
      RECT 4.650000  1.035000 4.970000 1.995000 ;
      RECT 5.140000  0.535000 5.310000 0.995000 ;
      RECT 5.140000  0.995000 6.015000 1.325000 ;
      RECT 5.140000  1.325000 5.310000 2.165000 ;
      RECT 5.480000  1.530000 6.375000 1.905000 ;
      RECT 5.490000  2.135000 5.805000 2.635000 ;
      RECT 5.585000  0.085000 5.795000 0.615000 ;
      RECT 6.035000  1.905000 6.375000 2.465000 ;
      RECT 6.055000  0.300000 6.385000 0.825000 ;
      RECT 6.185000  0.825000 6.385000 0.995000 ;
      RECT 6.185000  0.995000 6.935000 1.325000 ;
      RECT 6.185000  1.325000 6.375000 1.530000 ;
      RECT 6.545000  1.625000 6.715000 2.635000 ;
      RECT 6.555000  0.085000 6.725000 0.695000 ;
      RECT 7.385000  1.720000 7.555000 2.635000 ;
      RECT 7.395000  0.085000 7.565000 0.600000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.630000  1.785000 0.800000 1.955000 ;
      RECT 1.025000  1.445000 1.195000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.215000  1.445000 2.385000 1.615000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.730000  1.785000 2.900000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.300000  1.785000 4.470000 1.955000 ;
      RECT 4.735000  1.445000 4.905000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 0.570000 1.755000 0.860000 1.800000 ;
      RECT 0.570000 1.800000 4.530000 1.940000 ;
      RECT 0.570000 1.940000 0.860000 1.985000 ;
      RECT 0.965000 1.415000 1.255000 1.460000 ;
      RECT 0.965000 1.460000 4.965000 1.600000 ;
      RECT 0.965000 1.600000 1.255000 1.645000 ;
      RECT 2.155000 1.415000 2.445000 1.460000 ;
      RECT 2.155000 1.600000 2.445000 1.645000 ;
      RECT 2.670000 1.755000 2.960000 1.800000 ;
      RECT 2.670000 1.940000 2.960000 1.985000 ;
      RECT 4.240000 1.755000 4.530000 1.800000 ;
      RECT 4.240000 1.940000 4.530000 1.985000 ;
      RECT 4.675000 1.415000 4.965000 1.460000 ;
      RECT 4.675000 1.600000 4.965000 1.645000 ;
  END
END sky130_fd_sc_hd__dfxtp_2
MACRO sky130_fd_sc_hd__decap_3
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_3 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.085000  0.085000 1.295000 0.835000 ;
      RECT 0.085000  0.835000 0.605000 1.375000 ;
      RECT 0.085000  1.545000 1.295000 2.635000 ;
      RECT 0.775000  1.005000 1.295000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_3
MACRO sky130_fd_sc_hd__decap_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.085000 1.755000 0.855000 ;
      RECT 0.085000  0.855000 0.835000 1.375000 ;
      RECT 0.085000  1.545000 1.755000 2.635000 ;
      RECT 1.005000  1.025000 1.755000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_4
MACRO sky130_fd_sc_hd__decap_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.085000 2.675000 0.855000 ;
      RECT 0.085000  0.855000 1.295000 1.375000 ;
      RECT 0.085000  1.545000 2.675000 2.635000 ;
      RECT 1.465000  1.025000 2.675000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_6
MACRO sky130_fd_sc_hd__decap_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.085000 5.430000 0.855000 ;
      RECT 0.085000  0.855000 2.665000 1.375000 ;
      RECT 0.085000  1.545000 5.430000 2.635000 ;
      RECT 2.835000  1.025000 5.430000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_12
MACRO sky130_fd_sc_hd__decap_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__decap_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 3.595000 0.855000 ;
      RECT 0.085000  0.855000 1.735000 1.375000 ;
      RECT 0.085000  1.545000 3.595000 2.635000 ;
      RECT 1.905000  1.025000 3.595000 1.545000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__decap_8
MACRO sky130_fd_sc_hd__a21o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.660000 1.015000 2.185000 1.325000 ;
        RECT 1.955000 0.375000 2.185000 1.015000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365000 0.995000 2.665000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 1.015000 1.480000 1.325000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.265000 0.355000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.525000  1.905000 0.865000 2.635000 ;
      RECT 0.545000  0.635000 1.775000 0.835000 ;
      RECT 0.545000  0.835000 0.835000 1.505000 ;
      RECT 0.545000  1.505000 1.315000 1.725000 ;
      RECT 0.615000  0.085000 1.285000 0.455000 ;
      RECT 1.045000  1.725000 1.315000 2.455000 ;
      RECT 1.465000  0.265000 1.775000 0.635000 ;
      RECT 1.495000  1.505000 2.655000 1.745000 ;
      RECT 1.495000  1.745000 1.725000 2.455000 ;
      RECT 1.895000  1.925000 2.225000 2.635000 ;
      RECT 2.365000  0.085000 2.655000 0.815000 ;
      RECT 2.395000  1.745000 2.655000 2.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__a21o_1
MACRO sky130_fd_sc_hd__a21o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.990000 1.010000 4.515000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.425000 1.010000 3.820000 1.275000 ;
        RECT 3.645000 1.275000 3.820000 1.510000 ;
        RECT 3.645000 1.510000 4.935000 1.680000 ;
        RECT 4.685000 1.055000 5.100000 1.290000 ;
        RECT 4.685000 1.290000 4.935000 1.510000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.395000 0.995000 2.705000 1.525000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.615000 1.735000 0.785000 ;
        RECT 0.145000 0.785000 0.630000 1.585000 ;
        RECT 0.145000 1.585000 1.735000 1.755000 ;
        RECT 0.625000 1.755000 0.795000 2.185000 ;
        RECT 1.485000 1.755000 1.735000 2.185000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.105000  0.085000 0.445000 0.445000 ;
      RECT 0.115000  1.935000 0.445000 2.635000 ;
      RECT 0.800000  0.995000 2.205000 1.325000 ;
      RECT 0.975000  0.085000 1.305000 0.445000 ;
      RECT 0.975000  1.935000 1.305000 2.635000 ;
      RECT 1.910000  0.085000 2.685000 0.445000 ;
      RECT 1.915000  1.515000 2.165000 2.635000 ;
      RECT 2.035000  0.615000 3.045000 0.670000 ;
      RECT 2.035000  0.670000 4.365000 0.785000 ;
      RECT 2.035000  0.785000 2.205000 0.995000 ;
      RECT 2.455000  1.695000 2.625000 2.295000 ;
      RECT 2.455000  2.295000 3.465000 2.465000 ;
      RECT 2.875000  0.255000 3.045000 0.615000 ;
      RECT 2.875000  0.785000 4.365000 0.840000 ;
      RECT 2.875000  0.840000 3.045000 2.125000 ;
      RECT 3.255000  0.085000 3.585000 0.445000 ;
      RECT 3.285000  1.445000 3.465000 1.850000 ;
      RECT 3.285000  1.850000 5.360000 2.020000 ;
      RECT 3.285000  2.020000 3.465000 2.295000 ;
      RECT 3.635000  2.275000 3.965000 2.635000 ;
      RECT 4.085000  0.405000 4.365000 0.670000 ;
      RECT 4.135000  2.020000 4.305000 2.465000 ;
      RECT 4.475000  2.275000 4.805000 2.635000 ;
      RECT 4.945000  0.085000 5.225000 0.885000 ;
      RECT 5.030000  2.020000 5.360000 2.395000 ;
      RECT 5.105000  1.460000 5.360000 1.850000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__a21o_4
MACRO sky130_fd_sc_hd__a21o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.240000 0.365000 2.620000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.810000 0.750000 3.125000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.995000 1.790000 1.410000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.635000 0.955000 0.825000 ;
        RECT 0.555000 0.825000 0.785000 2.465000 ;
        RECT 0.765000 0.255000 0.955000 0.635000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.095000  1.665000 0.385000 2.635000 ;
      RECT 0.265000  0.085000 0.595000 0.465000 ;
      RECT 0.955000  0.995000 1.295000 1.690000 ;
      RECT 0.955000  1.690000 1.790000 1.920000 ;
      RECT 0.955000  2.220000 1.285000 2.635000 ;
      RECT 1.125000  0.085000 1.455000 0.445000 ;
      RECT 1.125000  0.655000 1.865000 0.825000 ;
      RECT 1.125000  0.825000 1.295000 0.995000 ;
      RECT 1.475000  1.920000 1.790000 2.465000 ;
      RECT 1.675000  0.255000 1.865000 0.655000 ;
      RECT 1.960000  1.670000 3.075000 1.935000 ;
      RECT 1.960000  1.935000 2.185000 2.465000 ;
      RECT 2.355000  2.125000 2.685000 2.635000 ;
      RECT 2.805000  0.085000 3.135000 0.565000 ;
      RECT 2.855000  1.935000 3.075000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a21o_2
MACRO sky130_fd_sc_hd__or3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 2.350000 1.325000 ;
        RECT 1.525000 1.325000 1.770000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 2.125000 2.200000 2.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.325000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.860000 0.415000 3.135000 0.760000 ;
        RECT 2.860000 1.495000 3.135000 2.465000 ;
        RECT 2.965000 0.760000 3.135000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.905000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.515000  0.485000 0.845000 0.905000 ;
      RECT 0.595000  0.905000 0.845000 0.995000 ;
      RECT 0.595000  0.995000 1.310000 1.325000 ;
      RECT 0.595000  1.325000 0.765000 1.885000 ;
      RECT 1.025000  0.255000 1.285000 0.655000 ;
      RECT 1.025000  0.655000 2.690000 0.825000 ;
      RECT 1.025000  1.495000 1.355000 1.785000 ;
      RECT 1.025000  1.785000 2.200000 1.955000 ;
      RECT 1.455000  0.085000 1.785000 0.485000 ;
      RECT 1.955000  0.305000 2.125000 0.655000 ;
      RECT 2.030000  1.495000 2.690000 1.665000 ;
      RECT 2.030000  1.665000 2.200000 1.785000 ;
      RECT 2.295000  0.085000 2.670000 0.485000 ;
      RECT 2.370000  1.835000 2.650000 2.635000 ;
      RECT 2.520000  0.825000 2.690000 0.995000 ;
      RECT 2.520000  0.995000 2.795000 1.325000 ;
      RECT 2.520000  1.325000 2.690000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__or3b_1
MACRO sky130_fd_sc_hd__or3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 1.075000 2.230000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 2.125000 3.135000 2.365000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.640000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 0.265000 1.285000 0.595000 ;
        RECT 0.935000 0.595000 1.105000 1.495000 ;
        RECT 0.935000 1.495000 1.330000 1.700000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.290000 0.345000 0.735000 ;
      RECT 0.085000  0.735000 0.765000 0.905000 ;
      RECT 0.085000  1.810000 0.765000 1.870000 ;
      RECT 0.085000  1.870000 2.660000 1.955000 ;
      RECT 0.085000  1.955000 1.720000 2.040000 ;
      RECT 0.085000  2.040000 0.345000 2.220000 ;
      RECT 0.550000  2.210000 0.910000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.565000 ;
      RECT 0.595000  0.905000 0.765000 1.810000 ;
      RECT 1.275000  0.765000 3.135000 0.825000 ;
      RECT 1.275000  0.825000 2.160000 0.905000 ;
      RECT 1.275000  0.905000 1.595000 0.935000 ;
      RECT 1.275000  0.935000 1.445000 1.325000 ;
      RECT 1.425000  0.735000 3.135000 0.765000 ;
      RECT 1.425000  2.210000 1.755000 2.635000 ;
      RECT 1.520000  0.085000 1.690000 0.565000 ;
      RECT 1.550000  1.785000 2.660000 1.870000 ;
      RECT 1.990000  0.305000 2.160000 0.655000 ;
      RECT 1.990000  0.655000 3.135000 0.735000 ;
      RECT 2.330000  0.085000 2.660000 0.485000 ;
      RECT 2.490000  0.995000 2.790000 1.325000 ;
      RECT 2.490000  1.325000 2.660000 1.785000 ;
      RECT 2.830000  0.305000 3.085000 0.605000 ;
      RECT 2.830000  0.605000 3.135000 0.655000 ;
      RECT 2.830000  1.495000 3.135000 1.925000 ;
      RECT 2.965000  0.825000 3.135000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__or3b_2
MACRO sky130_fd_sc_hd__or3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.400000 1.415000 2.720000 1.700000 ;
        RECT 2.535000 0.995000 2.720000 1.415000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.890000 0.995000 3.200000 1.700000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.640000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 0.735000 2.025000 0.905000 ;
        RECT 0.935000 0.905000 1.105000 1.415000 ;
        RECT 0.935000 1.415000 2.220000 1.700000 ;
        RECT 1.000000 0.285000 1.330000 0.735000 ;
        RECT 1.855000 0.255000 2.090000 0.585000 ;
        RECT 1.855000 0.585000 2.025000 0.735000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.290000 0.345000 0.735000 ;
      RECT 0.085000  0.735000 0.765000 0.905000 ;
      RECT 0.085000  1.810000 0.765000 1.870000 ;
      RECT 0.085000  1.870000 3.620000 2.040000 ;
      RECT 0.085000  2.040000 0.345000 2.220000 ;
      RECT 0.550000  2.210000 0.910000 2.635000 ;
      RECT 0.595000  0.905000 0.765000 1.810000 ;
      RECT 0.620000  0.085000 0.790000 0.565000 ;
      RECT 1.275000  1.075000 2.365000 1.245000 ;
      RECT 1.420000  2.210000 1.750000 2.635000 ;
      RECT 1.500000  0.085000 1.670000 0.565000 ;
      RECT 2.195000  0.720000 4.055000 0.825000 ;
      RECT 2.195000  0.825000 2.400000 0.890000 ;
      RECT 2.195000  0.890000 2.365000 1.075000 ;
      RECT 2.250000  0.655000 4.055000 0.720000 ;
      RECT 2.255000  2.210000 2.595000 2.635000 ;
      RECT 2.260000  0.085000 2.590000 0.485000 ;
      RECT 2.760000  0.305000 2.930000 0.655000 ;
      RECT 3.100000  0.085000 3.490000 0.485000 ;
      RECT 3.390000  0.995000 3.680000 1.325000 ;
      RECT 3.390000  1.325000 3.620000 1.870000 ;
      RECT 3.520000  2.210000 4.055000 2.425000 ;
      RECT 3.660000  0.305000 3.915000 0.605000 ;
      RECT 3.660000  0.605000 4.055000 0.655000 ;
      RECT 3.850000  0.825000 4.055000 2.210000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__or3b_4
MACRO sky130_fd_sc_hd__inv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.320000 1.075000 0.650000 1.315000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.720000 0.255000 1.050000 0.885000 ;
        RECT 0.720000 1.485000 1.050000 2.465000 ;
        RECT 0.820000 0.885000 1.050000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.320000  0.085000 0.550000 0.905000 ;
      RECT 0.340000  1.495000 0.550000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_1
MACRO sky130_fd_sc_hd__inv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.680000 1.075000 3.535000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 4.055000 0.905000 ;
        RECT 0.085000 0.905000 0.430000 1.495000 ;
        RECT 0.085000 1.495000 4.055000 1.665000 ;
        RECT 0.680000 0.255000 1.010000 0.715000 ;
        RECT 0.680000 1.665000 1.010000 2.465000 ;
        RECT 1.520000 0.255000 1.850000 0.715000 ;
        RECT 1.520000 1.665000 1.850000 2.465000 ;
        RECT 2.360000 0.255000 2.690000 0.715000 ;
        RECT 2.360000 1.665000 2.690000 2.465000 ;
        RECT 3.200000 0.255000 3.530000 0.715000 ;
        RECT 3.200000 1.665000 3.530000 2.465000 ;
        RECT 3.735000 0.905000 4.055000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.255000  0.085000 0.510000 0.545000 ;
      RECT 0.255000  1.835000 0.510000 2.635000 ;
      RECT 1.180000  0.085000 1.350000 0.545000 ;
      RECT 1.180000  1.835000 1.350000 2.635000 ;
      RECT 2.020000  0.085000 2.190000 0.545000 ;
      RECT 2.020000  1.835000 2.190000 2.635000 ;
      RECT 2.860000  0.085000 3.030000 0.545000 ;
      RECT 2.860000  1.835000 3.030000 2.635000 ;
      RECT 3.700000  0.085000 4.005000 0.545000 ;
      RECT 3.700000  1.835000 4.000000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_8
MACRO sky130_fd_sc_hd__inv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.735000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 0.255000 0.895000 0.725000 ;
        RECT 0.565000 0.725000 2.170000 0.905000 ;
        RECT 0.565000 1.495000 2.170000 1.665000 ;
        RECT 0.565000 1.665000 0.895000 2.465000 ;
        RECT 1.405000 0.255000 1.735000 0.725000 ;
        RECT 1.405000 1.665000 2.170000 1.685000 ;
        RECT 1.405000 1.685000 1.735000 2.465000 ;
        RECT 1.905000 0.905000 2.170000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.130000  0.085000 0.395000 0.545000 ;
      RECT 0.130000  1.495000 0.395000 2.635000 ;
      RECT 1.065000  0.085000 1.235000 0.545000 ;
      RECT 1.065000  1.835000 1.235000 2.635000 ;
      RECT 1.905000  0.085000 2.155000 0.550000 ;
      RECT 1.905000  2.175000 2.115000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_4
MACRO sky130_fd_sc_hd__inv_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.970000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.680000 1.075000 5.270000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.673000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 5.895000 0.905000 ;
        RECT 0.085000 0.905000 0.510000 1.495000 ;
        RECT 0.085000 1.495000 5.895000 1.665000 ;
        RECT 0.680000 0.255000 1.010000 0.715000 ;
        RECT 0.680000 1.665000 1.010000 2.465000 ;
        RECT 1.520000 0.255000 1.850000 0.715000 ;
        RECT 1.520000 1.665000 1.850000 2.465000 ;
        RECT 2.360000 0.255000 2.690000 0.715000 ;
        RECT 2.360000 1.665000 2.690000 2.465000 ;
        RECT 3.200000 0.255000 3.530000 0.715000 ;
        RECT 3.200000 1.665000 3.530000 2.465000 ;
        RECT 4.040000 0.255000 4.370000 0.715000 ;
        RECT 4.040000 1.665000 4.370000 2.465000 ;
        RECT 4.880000 0.255000 5.210000 0.715000 ;
        RECT 4.880000 1.665000 5.210000 2.465000 ;
        RECT 5.545000 0.905000 5.895000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.255000  0.085000 0.510000 0.545000 ;
      RECT 0.255000  1.835000 0.510000 2.635000 ;
      RECT 1.180000  0.085000 1.350000 0.545000 ;
      RECT 1.180000  1.835000 1.350000 2.635000 ;
      RECT 2.020000  0.085000 2.190000 0.545000 ;
      RECT 2.020000  1.835000 2.190000 2.635000 ;
      RECT 2.860000  0.085000 3.030000 0.545000 ;
      RECT 2.860000  1.835000 3.030000 2.635000 ;
      RECT 3.700000  0.085000 3.870000 0.545000 ;
      RECT 3.700000  1.835000 3.870000 2.635000 ;
      RECT 4.540000  0.085000 4.710000 0.545000 ;
      RECT 4.540000  1.835000 4.710000 2.635000 ;
      RECT 5.555000  0.085000 5.895000 0.545000 ;
      RECT 5.555000  1.835000 5.895000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_12
MACRO sky130_fd_sc_hd__inv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  3.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 5.525000 1.315000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 0.255000 0.910000 0.715000 ;
        RECT 0.580000 0.715000 6.790000 0.905000 ;
        RECT 0.580000 1.495000 6.790000 1.665000 ;
        RECT 0.580000 1.665000 0.910000 2.465000 ;
        RECT 1.420000 0.255000 1.750000 0.715000 ;
        RECT 1.420000 1.665000 1.750000 2.465000 ;
        RECT 2.260000 0.255000 2.590000 0.715000 ;
        RECT 2.260000 1.665000 2.590000 2.465000 ;
        RECT 3.100000 0.255000 3.430000 0.715000 ;
        RECT 3.100000 1.665000 3.430000 2.465000 ;
        RECT 3.940000 0.255000 4.270000 0.715000 ;
        RECT 3.940000 1.665000 4.270000 2.465000 ;
        RECT 4.780000 0.255000 5.110000 0.715000 ;
        RECT 4.780000 1.665000 5.110000 2.465000 ;
        RECT 5.620000 0.255000 5.950000 0.715000 ;
        RECT 5.620000 1.665000 5.950000 2.465000 ;
        RECT 6.460000 0.255000 6.790000 0.715000 ;
        RECT 6.460000 0.905000 6.790000 1.495000 ;
        RECT 6.460000 1.665000 6.790000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.180000  0.085000 0.410000 0.885000 ;
      RECT 0.200000  1.485000 0.410000 2.635000 ;
      RECT 1.080000  0.085000 1.250000 0.545000 ;
      RECT 1.080000  1.835000 1.250000 2.635000 ;
      RECT 1.920000  0.085000 2.090000 0.545000 ;
      RECT 1.920000  1.835000 2.090000 2.635000 ;
      RECT 2.760000  0.085000 2.930000 0.545000 ;
      RECT 2.760000  1.835000 2.930000 2.635000 ;
      RECT 3.600000  0.085000 3.770000 0.545000 ;
      RECT 3.600000  1.835000 3.770000 2.635000 ;
      RECT 4.440000  0.085000 4.610000 0.545000 ;
      RECT 4.440000  1.835000 4.610000 2.635000 ;
      RECT 5.280000  0.085000 5.450000 0.545000 ;
      RECT 5.280000  1.835000 5.450000 2.635000 ;
      RECT 6.120000  0.085000 6.290000 0.545000 ;
      RECT 6.120000  1.835000 6.290000 2.635000 ;
      RECT 6.960000  0.085000 7.170000 0.885000 ;
      RECT 6.960000  1.835000 7.170000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_16
MACRO sky130_fd_sc_hd__inv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 0.435000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 0.255000 0.855000 0.885000 ;
        RECT 0.525000 1.485000 0.855000 2.465000 ;
        RECT 0.605000 0.885000 0.855000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.125000  0.085000 0.355000 0.905000 ;
      RECT 0.125000  1.495000 0.355000 2.635000 ;
      RECT 1.025000  0.085000 1.235000 0.905000 ;
      RECT 1.025000  1.495000 1.235000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_2
MACRO sky130_fd_sc_hd__inv_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.485000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 2.615000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.336500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.685000 1.495000 3.135000 1.665000 ;
        RECT 0.685000 1.665000 1.015000 2.465000 ;
        RECT 0.765000 0.255000 0.935000 0.725000 ;
        RECT 0.765000 0.725000 3.135000 0.905000 ;
        RECT 1.525000 1.665000 1.855000 2.465000 ;
        RECT 1.605000 0.255000 1.775000 0.725000 ;
        RECT 2.365000 1.665000 3.135000 1.685000 ;
        RECT 2.365000 1.685000 2.695000 2.465000 ;
        RECT 2.445000 0.255000 2.615000 0.725000 ;
        RECT 2.785000 0.905000 3.135000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.130000  0.085000 0.395000 0.545000 ;
      RECT 0.130000  1.495000 0.425000 2.635000 ;
      RECT 1.185000  0.085000 1.355000 0.545000 ;
      RECT 1.185000  1.835000 1.355000 2.635000 ;
      RECT 2.025000  0.085000 2.195000 0.545000 ;
      RECT 2.025000  1.835000 2.195000 2.635000 ;
      RECT 2.785000  0.085000 3.035000 0.550000 ;
      RECT 2.865000  2.175000 3.035000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__inv_6
MACRO sky130_fd_sc_hd__dfrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855000 0.265000 9.110000 0.795000 ;
        RECT 8.855000 1.445000 9.110000 2.325000 ;
        RECT 8.900000 0.795000 9.110000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.090000  0.345000 0.345000 0.635000 ;
      RECT 0.090000  0.635000 0.840000 0.805000 ;
      RECT 0.090000  1.795000 0.840000 1.965000 ;
      RECT 0.090000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 2.465000 ;
      RECT 1.545000  0.085000 1.875000 0.445000 ;
      RECT 1.850000  2.175000 2.100000 2.635000 ;
      RECT 2.045000  0.305000 2.540000 0.475000 ;
      RECT 2.045000  0.475000 2.215000 1.835000 ;
      RECT 2.045000  1.835000 2.440000 2.005000 ;
      RECT 2.270000  2.005000 2.440000 2.135000 ;
      RECT 2.270000  2.135000 2.520000 2.465000 ;
      RECT 2.385000  0.765000 2.735000 1.385000 ;
      RECT 2.610000  1.575000 3.075000 1.965000 ;
      RECT 2.735000  2.135000 3.415000 2.465000 ;
      RECT 2.745000  0.305000 3.600000 0.475000 ;
      RECT 2.905000  0.765000 3.260000 0.985000 ;
      RECT 2.905000  0.985000 3.075000 1.575000 ;
      RECT 3.245000  1.185000 4.935000 1.355000 ;
      RECT 3.245000  1.355000 3.415000 2.135000 ;
      RECT 3.430000  0.475000 3.600000 1.185000 ;
      RECT 3.585000  1.865000 4.660000 2.035000 ;
      RECT 3.585000  2.035000 3.755000 2.375000 ;
      RECT 3.775000  1.525000 5.275000 1.695000 ;
      RECT 3.990000  2.205000 4.320000 2.635000 ;
      RECT 4.475000  0.085000 4.805000 0.545000 ;
      RECT 4.490000  2.035000 4.660000 2.375000 ;
      RECT 4.765000  1.005000 4.935000 1.185000 ;
      RECT 4.955000  2.175000 5.325000 2.635000 ;
      RECT 5.015000  0.275000 5.365000 0.445000 ;
      RECT 5.015000  0.445000 5.275000 0.835000 ;
      RECT 5.105000  0.835000 5.275000 1.525000 ;
      RECT 5.105000  1.695000 5.275000 1.835000 ;
      RECT 5.105000  1.835000 5.665000 2.005000 ;
      RECT 5.465000  0.705000 5.675000 1.495000 ;
      RECT 5.465000  1.495000 6.140000 1.655000 ;
      RECT 5.465000  1.655000 6.430000 1.665000 ;
      RECT 5.495000  2.005000 5.665000 2.465000 ;
      RECT 5.585000  0.255000 6.535000 0.535000 ;
      RECT 5.845000  0.705000 6.195000 1.325000 ;
      RECT 5.900000  2.125000 6.770000 2.465000 ;
      RECT 5.970000  1.665000 6.430000 1.955000 ;
      RECT 6.365000  0.535000 6.535000 1.315000 ;
      RECT 6.365000  1.315000 6.770000 1.485000 ;
      RECT 6.600000  1.485000 6.770000 1.575000 ;
      RECT 6.600000  1.575000 7.820000 1.745000 ;
      RECT 6.600000  1.745000 6.770000 2.125000 ;
      RECT 6.705000  0.085000 6.895000 0.525000 ;
      RECT 6.705000  0.695000 7.235000 0.865000 ;
      RECT 6.705000  0.865000 6.925000 1.145000 ;
      RECT 6.940000  2.175000 7.190000 2.635000 ;
      RECT 7.065000  0.295000 8.135000 0.465000 ;
      RECT 7.065000  0.465000 7.235000 0.695000 ;
      RECT 7.360000  1.915000 8.160000 2.085000 ;
      RECT 7.360000  2.085000 7.530000 2.375000 ;
      RECT 7.710000  2.255000 8.040000 2.635000 ;
      RECT 7.815000  0.465000 8.135000 0.820000 ;
      RECT 7.815000  0.820000 8.140000 0.995000 ;
      RECT 7.815000  0.995000 8.730000 1.295000 ;
      RECT 7.990000  1.295000 8.730000 1.325000 ;
      RECT 7.990000  1.325000 8.160000 1.915000 ;
      RECT 8.380000  0.085000 8.685000 0.545000 ;
      RECT 8.380000  1.495000 8.685000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.655000  1.785000 0.825000 1.955000 ;
      RECT 1.015000  1.105000 1.185000 1.275000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.105000 2.615000 1.275000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  1.785000 3.075000 1.955000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.025000  1.105000 6.195000 1.275000 ;
      RECT 6.025000  1.785000 6.195000 1.955000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 0.595000 1.755000 0.885000 1.800000 ;
      RECT 0.595000 1.800000 6.255000 1.940000 ;
      RECT 0.595000 1.940000 0.885000 1.985000 ;
      RECT 0.955000 1.075000 1.245000 1.120000 ;
      RECT 0.955000 1.120000 6.255000 1.260000 ;
      RECT 0.955000 1.260000 1.245000 1.305000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrtn_1
MACRO sky130_fd_sc_hd__sdfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.88000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.140000 0.265000 11.400000 0.795000 ;
        RECT 11.140000 1.460000 11.400000 2.325000 ;
        RECT 11.150000 1.445000 11.400000 1.460000 ;
        RECT 11.190000 0.795000 11.400000 0.995000 ;
        RECT 11.190000 0.995000 12.240000 1.325000 ;
        RECT 11.190000 1.325000 11.400000 1.445000 ;
        RECT 11.990000 0.265000 12.240000 0.995000 ;
        RECT 11.990000 1.325000 12.240000 2.325000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
      LAYER mcon ;
        RECT 6.865000 0.765000 7.035000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
      LAYER mcon ;
        RECT 9.690000 1.105000  9.860000 1.275000 ;
        RECT 9.945000 0.765000 10.115000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.880000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215000 -0.010000 0.235000 0.015000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  1.970000 1.425000 ;
        RECT -0.190000 1.425000 13.070000 2.910000 ;
        RECT  4.405000 1.305000 13.070000 1.425000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.880000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.880000 0.085000 ;
      RECT  0.000000  2.635000 12.880000 2.805000 ;
      RECT  0.090000  1.795000  0.865000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.530000  2.135000  0.860000 2.635000 ;
      RECT  0.660000  0.805000  0.835000 0.995000 ;
      RECT  0.660000  0.995000  0.975000 1.325000 ;
      RECT  0.660000  1.325000  0.865000 1.795000 ;
      RECT  1.015000  0.345000  1.315000 0.675000 ;
      RECT  1.035000  1.730000  1.315000 1.900000 ;
      RECT  1.035000  1.900000  1.205000 2.465000 ;
      RECT  1.145000  0.675000  1.315000 1.730000 ;
      RECT  1.535000  0.395000  1.705000 0.730000 ;
      RECT  1.535000  0.730000  2.225000 0.900000 ;
      RECT  1.875000  0.085000  2.205000 0.560000 ;
      RECT  1.900000  2.055000  2.150000 2.400000 ;
      RECT  1.980000  1.260000  2.470000 1.455000 ;
      RECT  1.980000  1.455000  2.150000 2.055000 ;
      RECT  2.055000  0.900000  2.225000 0.995000 ;
      RECT  2.055000  0.995000  3.085000 1.185000 ;
      RECT  2.055000  1.185000  2.470000 1.260000 ;
      RECT  2.320000  2.040000  2.490000 2.635000 ;
      RECT  2.395000  0.085000  2.725000 0.825000 ;
      RECT  2.915000  0.255000  3.850000 0.425000 ;
      RECT  2.915000  0.425000  3.085000 0.995000 ;
      RECT  3.255000  0.675000  3.425000 1.015000 ;
      RECT  3.255000  1.015000  3.460000 1.185000 ;
      RECT  3.290000  1.185000  3.460000 1.935000 ;
      RECT  3.290000  1.935000  5.075000 2.105000 ;
      RECT  3.460000  2.105000  3.630000 2.465000 ;
      RECT  3.680000  0.425000  3.850000 1.685000 ;
      RECT  4.300000  2.275000  4.630000 2.635000 ;
      RECT  4.445000  0.085000  4.775000 0.540000 ;
      RECT  4.565000  0.715000  5.145000 0.895000 ;
      RECT  4.565000  0.895000  4.735000 1.935000 ;
      RECT  4.905000  1.065000  5.075000 1.395000 ;
      RECT  4.905000  2.105000  5.075000 2.185000 ;
      RECT  4.905000  2.185000  5.275000 2.435000 ;
      RECT  4.975000  0.335000  5.315000 0.505000 ;
      RECT  4.975000  0.505000  5.145000 0.715000 ;
      RECT  5.245000  1.575000  5.495000 1.955000 ;
      RECT  5.325000  0.705000  5.975000 1.035000 ;
      RECT  5.325000  1.035000  5.495000 1.575000 ;
      RECT  5.470000  2.135000  5.835000 2.465000 ;
      RECT  5.485000  0.305000  6.335000 0.475000 ;
      RECT  5.665000  1.215000  7.375000 1.385000 ;
      RECT  5.665000  1.385000  5.835000 2.135000 ;
      RECT  6.005000  1.935000  7.165000 2.105000 ;
      RECT  6.005000  2.105000  6.175000 2.375000 ;
      RECT  6.165000  0.475000  6.335000 1.215000 ;
      RECT  6.285000  1.595000  7.715000 1.765000 ;
      RECT  6.410000  2.355000  6.740000 2.635000 ;
      RECT  6.915000  0.085000  7.245000 0.545000 ;
      RECT  6.995000  2.105000  7.165000 2.375000 ;
      RECT  7.205000  1.005000  7.375000 1.215000 ;
      RECT  7.375000  2.175000  7.745000 2.635000 ;
      RECT  7.455000  0.275000  7.785000 0.445000 ;
      RECT  7.455000  0.445000  7.715000 0.835000 ;
      RECT  7.455000  1.765000  7.715000 1.835000 ;
      RECT  7.455000  1.835000  8.140000 2.005000 ;
      RECT  7.545000  0.835000  7.715000 1.595000 ;
      RECT  7.885000  0.705000  8.095000 1.495000 ;
      RECT  7.885000  1.495000  8.520000 1.655000 ;
      RECT  7.885000  1.655000  8.870000 1.665000 ;
      RECT  7.970000  2.005000  8.140000 2.465000 ;
      RECT  8.005000  0.255000  8.915000 0.535000 ;
      RECT  8.310000  1.665000  8.870000 1.935000 ;
      RECT  8.310000  1.935000  8.840000 1.955000 ;
      RECT  8.320000  2.125000  9.190000 2.465000 ;
      RECT  8.405000  0.920000  8.575000 1.325000 ;
      RECT  8.745000  0.535000  8.915000 1.315000 ;
      RECT  8.745000  1.315000  9.210000 1.485000 ;
      RECT  9.015000  2.035000  9.210000 2.115000 ;
      RECT  9.015000  2.115000  9.190000 2.125000 ;
      RECT  9.040000  1.485000  9.210000 1.575000 ;
      RECT  9.040000  1.575000 10.205000 1.745000 ;
      RECT  9.040000  1.745000  9.210000 2.035000 ;
      RECT  9.085000  0.085000  9.255000 0.525000 ;
      RECT  9.125000  0.695000  9.655000 0.865000 ;
      RECT  9.125000  0.865000  9.295000 1.145000 ;
      RECT  9.360000  2.195000  9.610000 2.635000 ;
      RECT  9.485000  0.295000 10.515000 0.465000 ;
      RECT  9.485000  0.465000  9.655000 0.695000 ;
      RECT  9.780000  1.915000 10.545000 2.085000 ;
      RECT  9.780000  2.085000  9.950000 2.375000 ;
      RECT 10.120000  2.255000 10.450000 2.635000 ;
      RECT 10.345000  0.465000 10.515000 0.995000 ;
      RECT 10.345000  0.995000 11.020000 1.295000 ;
      RECT 10.375000  1.295000 11.020000 1.325000 ;
      RECT 10.375000  1.325000 10.545000 1.915000 ;
      RECT 10.720000  0.085000 10.890000 0.545000 ;
      RECT 10.720000  1.495000 10.970000 2.635000 ;
      RECT 11.570000  0.085000 11.740000 0.545000 ;
      RECT 11.570000  1.495000 11.820000 2.635000 ;
      RECT 12.410000  0.085000 12.580000 0.545000 ;
      RECT 12.410000  1.495000 12.660000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.805000  1.105000  0.975000 1.275000 ;
      RECT  1.035000  1.785000  1.205000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.905000  1.105000  5.075000 1.275000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.325000  1.785000  5.495000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.405000  1.105000  8.575000 1.275000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.445000  1.785000  8.615000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
    LAYER met1 ;
      RECT 0.745000 1.075000 1.035000 1.120000 ;
      RECT 0.745000 1.120000 8.635000 1.260000 ;
      RECT 0.745000 1.260000 1.035000 1.305000 ;
      RECT 0.970000 1.755000 1.270000 1.800000 ;
      RECT 0.970000 1.800000 8.675000 1.940000 ;
      RECT 0.970000 1.940000 1.270000 1.985000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrtp_4
MACRO sky130_fd_sc_hd__sdfrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.140000 0.265000 11.400000 0.795000 ;
        RECT 11.140000 1.460000 11.400000 2.325000 ;
        RECT 11.150000 1.445000 11.400000 1.460000 ;
        RECT 11.190000 0.795000 11.400000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
      LAYER mcon ;
        RECT 6.865000 0.765000 7.035000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
      LAYER mcon ;
        RECT 9.690000 1.105000  9.860000 1.275000 ;
        RECT 9.945000 0.765000 10.115000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215000 -0.010000 0.235000 0.015000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  1.970000 1.425000 ;
        RECT -0.190000 1.425000 12.150000 2.910000 ;
        RECT  4.405000 1.305000 12.150000 1.425000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.090000  1.795000  0.865000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.530000  2.135000  0.860000 2.635000 ;
      RECT  0.660000  0.805000  0.835000 0.995000 ;
      RECT  0.660000  0.995000  0.975000 1.325000 ;
      RECT  0.660000  1.325000  0.865000 1.795000 ;
      RECT  1.015000  0.345000  1.315000 0.675000 ;
      RECT  1.035000  1.730000  1.315000 1.900000 ;
      RECT  1.035000  1.900000  1.205000 2.465000 ;
      RECT  1.145000  0.675000  1.315000 1.730000 ;
      RECT  1.535000  0.395000  1.705000 0.730000 ;
      RECT  1.535000  0.730000  2.225000 0.900000 ;
      RECT  1.875000  0.085000  2.205000 0.560000 ;
      RECT  1.900000  2.055000  2.150000 2.400000 ;
      RECT  1.980000  1.260000  2.470000 1.455000 ;
      RECT  1.980000  1.455000  2.150000 2.055000 ;
      RECT  2.055000  0.900000  2.225000 0.995000 ;
      RECT  2.055000  0.995000  3.085000 1.185000 ;
      RECT  2.055000  1.185000  2.470000 1.260000 ;
      RECT  2.320000  2.040000  2.490000 2.635000 ;
      RECT  2.395000  0.085000  2.725000 0.825000 ;
      RECT  2.915000  0.255000  3.850000 0.425000 ;
      RECT  2.915000  0.425000  3.085000 0.995000 ;
      RECT  3.255000  0.675000  3.425000 1.015000 ;
      RECT  3.255000  1.015000  3.460000 1.185000 ;
      RECT  3.290000  1.185000  3.460000 1.935000 ;
      RECT  3.290000  1.935000  5.075000 2.105000 ;
      RECT  3.460000  2.105000  3.630000 2.465000 ;
      RECT  3.680000  0.425000  3.850000 1.685000 ;
      RECT  4.300000  2.275000  4.630000 2.635000 ;
      RECT  4.445000  0.085000  4.775000 0.540000 ;
      RECT  4.565000  0.715000  5.145000 0.895000 ;
      RECT  4.565000  0.895000  4.735000 1.935000 ;
      RECT  4.905000  1.065000  5.075000 1.395000 ;
      RECT  4.905000  2.105000  5.075000 2.185000 ;
      RECT  4.905000  2.185000  5.275000 2.435000 ;
      RECT  4.975000  0.335000  5.315000 0.505000 ;
      RECT  4.975000  0.505000  5.145000 0.715000 ;
      RECT  5.245000  1.575000  5.495000 1.955000 ;
      RECT  5.325000  0.705000  5.975000 1.035000 ;
      RECT  5.325000  1.035000  5.495000 1.575000 ;
      RECT  5.470000  2.135000  5.835000 2.465000 ;
      RECT  5.485000  0.305000  6.335000 0.475000 ;
      RECT  5.665000  1.215000  7.375000 1.385000 ;
      RECT  5.665000  1.385000  5.835000 2.135000 ;
      RECT  6.005000  1.935000  7.165000 2.105000 ;
      RECT  6.005000  2.105000  6.175000 2.375000 ;
      RECT  6.165000  0.475000  6.335000 1.215000 ;
      RECT  6.285000  1.595000  7.715000 1.765000 ;
      RECT  6.410000  2.355000  6.740000 2.635000 ;
      RECT  6.915000  0.085000  7.245000 0.545000 ;
      RECT  6.995000  2.105000  7.165000 2.375000 ;
      RECT  7.205000  1.005000  7.375000 1.215000 ;
      RECT  7.375000  2.175000  7.745000 2.635000 ;
      RECT  7.455000  0.275000  7.785000 0.445000 ;
      RECT  7.455000  0.445000  7.715000 0.835000 ;
      RECT  7.455000  1.765000  7.715000 1.835000 ;
      RECT  7.455000  1.835000  8.140000 2.005000 ;
      RECT  7.545000  0.835000  7.715000 1.595000 ;
      RECT  7.885000  0.705000  8.095000 1.495000 ;
      RECT  7.885000  1.495000  8.520000 1.655000 ;
      RECT  7.885000  1.655000  8.870000 1.665000 ;
      RECT  7.970000  2.005000  8.140000 2.465000 ;
      RECT  8.005000  0.255000  8.915000 0.535000 ;
      RECT  8.310000  1.665000  8.870000 1.935000 ;
      RECT  8.310000  1.935000  8.840000 1.955000 ;
      RECT  8.320000  2.125000  9.190000 2.465000 ;
      RECT  8.405000  0.920000  8.575000 1.325000 ;
      RECT  8.745000  0.535000  8.915000 1.315000 ;
      RECT  8.745000  1.315000  9.210000 1.485000 ;
      RECT  9.015000  2.035000  9.210000 2.115000 ;
      RECT  9.015000  2.115000  9.190000 2.125000 ;
      RECT  9.040000  1.485000  9.210000 1.575000 ;
      RECT  9.040000  1.575000 10.205000 1.745000 ;
      RECT  9.040000  1.745000  9.210000 2.035000 ;
      RECT  9.085000  0.085000  9.255000 0.525000 ;
      RECT  9.125000  0.695000  9.655000 0.865000 ;
      RECT  9.125000  0.865000  9.295000 1.145000 ;
      RECT  9.360000  2.195000  9.610000 2.635000 ;
      RECT  9.485000  0.295000 10.515000 0.465000 ;
      RECT  9.485000  0.465000  9.655000 0.695000 ;
      RECT  9.780000  1.915000 10.545000 2.085000 ;
      RECT  9.780000  2.085000  9.950000 2.375000 ;
      RECT 10.120000  2.255000 10.450000 2.635000 ;
      RECT 10.345000  0.465000 10.515000 0.995000 ;
      RECT 10.345000  0.995000 11.020000 1.295000 ;
      RECT 10.375000  1.295000 11.020000 1.325000 ;
      RECT 10.375000  1.325000 10.545000 1.915000 ;
      RECT 10.720000  0.085000 10.890000 0.545000 ;
      RECT 10.720000  1.495000 10.970000 2.635000 ;
      RECT 11.570000  0.085000 11.740000 0.545000 ;
      RECT 11.570000  1.495000 11.820000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.805000  1.105000  0.975000 1.275000 ;
      RECT  1.035000  1.785000  1.205000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.905000  1.105000  5.075000 1.275000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.325000  1.785000  5.495000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.405000  1.105000  8.575000 1.275000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.445000  1.785000  8.615000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.745000 1.075000 1.035000 1.120000 ;
      RECT 0.745000 1.120000 8.635000 1.260000 ;
      RECT 0.745000 1.260000 1.035000 1.305000 ;
      RECT 0.970000 1.755000 1.270000 1.800000 ;
      RECT 0.970000 1.800000 8.675000 1.940000 ;
      RECT 0.970000 1.940000 1.270000 1.985000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrtp_2
MACRO sky130_fd_sc_hd__sdfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.50000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.140000 0.265000 11.400000 0.795000 ;
        RECT 11.140000 1.460000 11.400000 2.325000 ;
        RECT 11.150000 1.445000 11.400000 1.460000 ;
        RECT 11.190000 0.795000 11.400000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
      LAYER mcon ;
        RECT 6.865000 0.765000 7.035000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
      LAYER mcon ;
        RECT 9.690000 1.105000  9.860000 1.275000 ;
        RECT 9.945000 0.765000 10.115000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.500000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215000 -0.010000 0.235000 0.015000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  1.970000 1.425000 ;
        RECT -0.190000 1.425000 11.690000 2.910000 ;
        RECT  4.405000 1.305000 11.690000 1.425000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.500000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.500000 0.085000 ;
      RECT  0.000000  2.635000 11.500000 2.805000 ;
      RECT  0.090000  1.795000  0.865000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.530000  2.135000  0.860000 2.635000 ;
      RECT  0.660000  0.805000  0.835000 0.995000 ;
      RECT  0.660000  0.995000  0.975000 1.325000 ;
      RECT  0.660000  1.325000  0.865000 1.795000 ;
      RECT  1.015000  0.345000  1.315000 0.675000 ;
      RECT  1.035000  1.730000  1.315000 1.900000 ;
      RECT  1.035000  1.900000  1.205000 2.465000 ;
      RECT  1.145000  0.675000  1.315000 1.730000 ;
      RECT  1.535000  0.395000  1.705000 0.730000 ;
      RECT  1.535000  0.730000  2.225000 0.900000 ;
      RECT  1.875000  0.085000  2.205000 0.560000 ;
      RECT  1.900000  2.055000  2.150000 2.400000 ;
      RECT  1.980000  1.260000  2.470000 1.455000 ;
      RECT  1.980000  1.455000  2.150000 2.055000 ;
      RECT  2.055000  0.900000  2.225000 0.995000 ;
      RECT  2.055000  0.995000  3.085000 1.185000 ;
      RECT  2.055000  1.185000  2.470000 1.260000 ;
      RECT  2.320000  2.040000  2.490000 2.635000 ;
      RECT  2.395000  0.085000  2.725000 0.825000 ;
      RECT  2.915000  0.255000  3.850000 0.425000 ;
      RECT  2.915000  0.425000  3.085000 0.995000 ;
      RECT  3.255000  0.675000  3.425000 1.015000 ;
      RECT  3.255000  1.015000  3.460000 1.185000 ;
      RECT  3.290000  1.185000  3.460000 1.935000 ;
      RECT  3.290000  1.935000  5.075000 2.105000 ;
      RECT  3.460000  2.105000  3.630000 2.465000 ;
      RECT  3.680000  0.425000  3.850000 1.685000 ;
      RECT  4.300000  2.275000  4.630000 2.635000 ;
      RECT  4.445000  0.085000  4.775000 0.540000 ;
      RECT  4.565000  0.715000  5.145000 0.895000 ;
      RECT  4.565000  0.895000  4.735000 1.935000 ;
      RECT  4.905000  1.065000  5.075000 1.395000 ;
      RECT  4.905000  2.105000  5.075000 2.185000 ;
      RECT  4.905000  2.185000  5.275000 2.435000 ;
      RECT  4.975000  0.335000  5.315000 0.505000 ;
      RECT  4.975000  0.505000  5.145000 0.715000 ;
      RECT  5.245000  1.575000  5.495000 1.955000 ;
      RECT  5.325000  0.705000  5.975000 1.035000 ;
      RECT  5.325000  1.035000  5.495000 1.575000 ;
      RECT  5.470000  2.135000  5.835000 2.465000 ;
      RECT  5.485000  0.305000  6.335000 0.475000 ;
      RECT  5.665000  1.215000  7.375000 1.385000 ;
      RECT  5.665000  1.385000  5.835000 2.135000 ;
      RECT  6.005000  1.935000  7.165000 2.105000 ;
      RECT  6.005000  2.105000  6.175000 2.375000 ;
      RECT  6.165000  0.475000  6.335000 1.215000 ;
      RECT  6.285000  1.595000  7.715000 1.765000 ;
      RECT  6.410000  2.355000  6.740000 2.635000 ;
      RECT  6.915000  0.085000  7.245000 0.545000 ;
      RECT  6.995000  2.105000  7.165000 2.375000 ;
      RECT  7.205000  1.005000  7.375000 1.215000 ;
      RECT  7.375000  2.175000  7.745000 2.635000 ;
      RECT  7.455000  0.275000  7.785000 0.445000 ;
      RECT  7.455000  0.445000  7.715000 0.835000 ;
      RECT  7.455000  1.765000  7.715000 1.835000 ;
      RECT  7.455000  1.835000  8.140000 2.005000 ;
      RECT  7.545000  0.835000  7.715000 1.595000 ;
      RECT  7.885000  0.705000  8.095000 1.495000 ;
      RECT  7.885000  1.495000  8.520000 1.655000 ;
      RECT  7.885000  1.655000  8.870000 1.665000 ;
      RECT  7.970000  2.005000  8.140000 2.465000 ;
      RECT  8.005000  0.255000  8.915000 0.535000 ;
      RECT  8.310000  1.665000  8.870000 1.935000 ;
      RECT  8.310000  1.935000  8.840000 1.955000 ;
      RECT  8.320000  2.125000  9.190000 2.465000 ;
      RECT  8.405000  0.920000  8.575000 1.325000 ;
      RECT  8.745000  0.535000  8.915000 1.315000 ;
      RECT  8.745000  1.315000  9.210000 1.485000 ;
      RECT  9.015000  2.035000  9.210000 2.115000 ;
      RECT  9.015000  2.115000  9.190000 2.125000 ;
      RECT  9.040000  1.485000  9.210000 1.575000 ;
      RECT  9.040000  1.575000 10.205000 1.745000 ;
      RECT  9.040000  1.745000  9.210000 2.035000 ;
      RECT  9.085000  0.085000  9.255000 0.525000 ;
      RECT  9.125000  0.695000  9.655000 0.865000 ;
      RECT  9.125000  0.865000  9.295000 1.145000 ;
      RECT  9.360000  2.195000  9.610000 2.635000 ;
      RECT  9.485000  0.295000 10.515000 0.465000 ;
      RECT  9.485000  0.465000  9.655000 0.695000 ;
      RECT  9.780000  1.915000 10.545000 2.085000 ;
      RECT  9.780000  2.085000  9.950000 2.375000 ;
      RECT 10.120000  2.255000 10.450000 2.635000 ;
      RECT 10.345000  0.465000 10.515000 0.995000 ;
      RECT 10.345000  0.995000 11.020000 1.295000 ;
      RECT 10.375000  1.295000 11.020000 1.325000 ;
      RECT 10.375000  1.325000 10.545000 1.915000 ;
      RECT 10.720000  0.085000 10.890000 0.545000 ;
      RECT 10.720000  1.495000 10.970000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.805000  1.105000  0.975000 1.275000 ;
      RECT  1.035000  1.785000  1.205000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.905000  1.105000  5.075000 1.275000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.325000  1.785000  5.495000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.405000  1.105000  8.575000 1.275000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.445000  1.785000  8.615000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
    LAYER met1 ;
      RECT 0.745000 1.075000 1.035000 1.120000 ;
      RECT 0.745000 1.120000 8.635000 1.260000 ;
      RECT 0.745000 1.260000 1.035000 1.305000 ;
      RECT 0.970000 1.755000 1.270000 1.800000 ;
      RECT 0.970000 1.800000 8.675000 1.940000 ;
      RECT 0.970000 1.940000 1.270000 1.985000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrtp_1
MACRO sky130_fd_sc_hd__bufinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufinv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.505000 1.275000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715000 0.260000 3.045000 0.735000 ;
        RECT 2.715000 0.735000 6.355000 0.905000 ;
        RECT 2.715000 1.445000 6.355000 1.615000 ;
        RECT 2.715000 1.615000 3.045000 2.465000 ;
        RECT 3.555000 0.260000 3.885000 0.735000 ;
        RECT 3.555000 1.615000 3.885000 2.465000 ;
        RECT 4.395000 0.260000 4.725000 0.735000 ;
        RECT 4.395000 1.615000 4.725000 2.465000 ;
        RECT 5.235000 0.260000 5.565000 0.735000 ;
        RECT 5.235000 1.615000 5.565000 2.465000 ;
        RECT 5.970000 0.905000 6.355000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.085000 0.345000 0.905000 ;
      RECT 0.175000  1.445000 0.345000 2.635000 ;
      RECT 0.515000  0.260000 0.845000 0.905000 ;
      RECT 0.515000  1.545000 0.845000 2.465000 ;
      RECT 0.675000  0.905000 0.845000 1.075000 ;
      RECT 0.675000  1.075000 2.205000 1.275000 ;
      RECT 0.675000  1.275000 0.845000 1.545000 ;
      RECT 1.035000  0.260000 1.365000 0.735000 ;
      RECT 1.035000  0.735000 2.545000 0.905000 ;
      RECT 1.035000  1.445000 2.545000 1.615000 ;
      RECT 1.035000  1.615000 1.365000 2.465000 ;
      RECT 1.535000  0.085000 1.705000 0.565000 ;
      RECT 1.535000  1.785000 1.705000 2.635000 ;
      RECT 1.875000  0.260000 2.205000 0.735000 ;
      RECT 1.875000  1.615000 2.205000 2.465000 ;
      RECT 2.375000  0.085000 2.545000 0.565000 ;
      RECT 2.375000  0.905000 2.545000 1.075000 ;
      RECT 2.375000  1.075000 5.760000 1.275000 ;
      RECT 2.375000  1.275000 2.545000 1.445000 ;
      RECT 2.375000  1.785000 2.545000 2.635000 ;
      RECT 3.215000  0.085000 3.385000 0.565000 ;
      RECT 3.215000  1.835000 3.385000 2.635000 ;
      RECT 4.055000  0.085000 4.225000 0.565000 ;
      RECT 4.055000  1.835000 4.225000 2.635000 ;
      RECT 4.895000  0.085000 5.065000 0.565000 ;
      RECT 4.895000  1.835000 5.065000 2.635000 ;
      RECT 5.735000  0.085000 5.905000 0.565000 ;
      RECT 5.735000  1.835000 5.905000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__bufinv_8
MACRO sky130_fd_sc_hd__bufinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufinv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.265000 1.275000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  4.295000 0.255000  4.545000 0.260000 ;
        RECT  4.295000 0.260000  4.625000 0.735000 ;
        RECT  4.295000 0.735000 10.955000 0.905000 ;
        RECT  4.295000 1.445000 10.955000 1.615000 ;
        RECT  4.295000 1.615000  4.625000 2.465000 ;
        RECT  5.135000 0.260000  5.465000 0.735000 ;
        RECT  5.135000 1.615000  5.465000 2.465000 ;
        RECT  5.215000 0.255000  5.385000 0.260000 ;
        RECT  5.975000 0.260000  6.305000 0.735000 ;
        RECT  5.975000 1.615000  6.305000 2.465000 ;
        RECT  6.055000 0.255000  6.225000 0.260000 ;
        RECT  6.815000 0.260000  7.145000 0.735000 ;
        RECT  6.815000 1.615000  7.145000 2.465000 ;
        RECT  7.655000 0.260000  7.985000 0.735000 ;
        RECT  7.655000 1.615000  7.985000 2.465000 ;
        RECT  8.495000 0.260000  8.825000 0.735000 ;
        RECT  8.495000 1.615000  8.825000 2.465000 ;
        RECT  9.335000 0.260000  9.665000 0.735000 ;
        RECT  9.335000 1.615000  9.665000 2.465000 ;
        RECT 10.175000 0.260000 10.505000 0.735000 ;
        RECT 10.175000 1.615000 10.505000 2.465000 ;
        RECT 10.680000 0.905000 10.955000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.095000  0.260000  0.425000 0.735000 ;
      RECT  0.095000  0.735000  1.605000 0.905000 ;
      RECT  0.095000  1.445000  1.605000 1.615000 ;
      RECT  0.095000  1.615000  0.425000 2.465000 ;
      RECT  0.595000  0.085000  0.765000 0.565000 ;
      RECT  0.595000  1.785000  0.765000 2.635000 ;
      RECT  0.935000  0.260000  1.265000 0.735000 ;
      RECT  0.935000  1.615000  1.265000 2.465000 ;
      RECT  1.435000  0.085000  1.605000 0.565000 ;
      RECT  1.435000  0.905000  1.605000 1.075000 ;
      RECT  1.435000  1.075000  3.745000 1.275000 ;
      RECT  1.435000  1.275000  1.605000 1.445000 ;
      RECT  1.435000  1.785000  1.605000 2.635000 ;
      RECT  1.775000  0.260000  2.105000 0.735000 ;
      RECT  1.775000  0.735000  4.125000 0.905000 ;
      RECT  1.775000  1.445000  4.125000 1.615000 ;
      RECT  1.775000  1.615000  2.105000 2.465000 ;
      RECT  2.275000  0.085000  2.445000 0.565000 ;
      RECT  2.275000  1.835000  2.445000 2.635000 ;
      RECT  2.615000  0.260000  2.945000 0.735000 ;
      RECT  2.615000  1.615000  2.945000 2.465000 ;
      RECT  3.115000  0.085000  3.285000 0.565000 ;
      RECT  3.115000  1.835000  3.285000 2.635000 ;
      RECT  3.455000  0.260000  3.785000 0.735000 ;
      RECT  3.455000  1.615000  3.785000 2.465000 ;
      RECT  3.950000  0.905000  4.125000 1.075000 ;
      RECT  3.950000  1.075000 10.510000 1.275000 ;
      RECT  3.950000  1.275000  4.125000 1.445000 ;
      RECT  3.955000  0.085000  4.125000 0.565000 ;
      RECT  3.955000  1.835000  4.125000 2.635000 ;
      RECT  4.795000  0.085000  4.965000 0.565000 ;
      RECT  4.795000  1.835000  4.965000 2.635000 ;
      RECT  5.635000  0.085000  5.805000 0.565000 ;
      RECT  5.635000  1.835000  5.805000 2.635000 ;
      RECT  6.475000  0.085000  6.645000 0.565000 ;
      RECT  6.475000  1.835000  6.645000 2.635000 ;
      RECT  7.315000  0.085000  7.485000 0.565000 ;
      RECT  7.315000  1.835000  7.485000 2.635000 ;
      RECT  8.155000  0.085000  8.325000 0.565000 ;
      RECT  8.155000  1.835000  8.325000 2.635000 ;
      RECT  8.995000  0.085000  9.165000 0.565000 ;
      RECT  8.995000  1.835000  9.165000 2.635000 ;
      RECT  9.835000  0.085000 10.005000 0.565000 ;
      RECT  9.835000  1.835000 10.005000 2.635000 ;
      RECT 10.675000  0.085000 10.845000 0.565000 ;
      RECT 10.675000  1.835000 10.845000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
  END
END sky130_fd_sc_hd__bufinv_16
MACRO sky130_fd_sc_hd__sdfrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.50000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.355000 3.120000 1.785000 ;
        RECT 2.865000 1.785000 3.120000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.140000 0.265000 11.400000 0.795000 ;
        RECT 11.140000 1.460000 11.400000 2.325000 ;
        RECT 11.150000 1.445000 11.400000 1.460000 ;
        RECT 11.190000 0.795000 11.400000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505000 0.765000 7.035000 1.045000 ;
      LAYER mcon ;
        RECT 6.865000 0.765000 7.035000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525000 1.065000 10.115000 1.275000 ;
        RECT 9.825000 0.635000 10.115000 1.065000 ;
      LAYER mcon ;
        RECT 9.690000 1.105000  9.860000 1.275000 ;
        RECT 9.945000 0.765000 10.115000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445000 0.735000  7.095000 0.780000 ;
        RECT 6.445000 0.780000 10.175000 0.920000 ;
        RECT 6.445000 0.920000  7.095000 0.965000 ;
        RECT 9.630000 0.920000 10.175000 0.965000 ;
        RECT 9.630000 0.965000  9.920000 1.305000 ;
        RECT 9.885000 0.735000 10.175000 0.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.020000 0.285000 4.275000 0.710000 ;
        RECT 4.020000 0.710000 4.395000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.985000 1.730000 2.465000 ;
        RECT 1.485000 1.070000 1.730000 1.985000 ;
    END
  END SCE
  PIN CLK_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.500000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.215000 -0.010000 0.235000 0.015000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  1.970000 1.425000 ;
        RECT -0.190000 1.425000 11.690000 2.910000 ;
        RECT  4.405000 1.305000 11.690000 1.425000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.500000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.500000 0.085000 ;
      RECT  0.000000  2.635000 11.500000 2.805000 ;
      RECT  0.090000  1.795000  0.865000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.530000  2.135000  0.860000 2.635000 ;
      RECT  0.660000  0.805000  0.835000 0.995000 ;
      RECT  0.660000  0.995000  0.975000 1.325000 ;
      RECT  0.660000  1.325000  0.865000 1.795000 ;
      RECT  1.015000  0.345000  1.315000 0.675000 ;
      RECT  1.035000  1.730000  1.315000 1.900000 ;
      RECT  1.035000  1.900000  1.205000 2.465000 ;
      RECT  1.145000  0.675000  1.315000 1.730000 ;
      RECT  1.535000  0.395000  1.705000 0.730000 ;
      RECT  1.535000  0.730000  2.225000 0.900000 ;
      RECT  1.875000  0.085000  2.205000 0.560000 ;
      RECT  1.900000  2.055000  2.150000 2.400000 ;
      RECT  1.980000  1.260000  2.470000 1.455000 ;
      RECT  1.980000  1.455000  2.150000 2.055000 ;
      RECT  2.055000  0.900000  2.225000 0.995000 ;
      RECT  2.055000  0.995000  3.085000 1.185000 ;
      RECT  2.055000  1.185000  2.470000 1.260000 ;
      RECT  2.320000  2.040000  2.490000 2.635000 ;
      RECT  2.395000  0.085000  2.725000 0.825000 ;
      RECT  2.915000  0.255000  3.850000 0.425000 ;
      RECT  2.915000  0.425000  3.085000 0.995000 ;
      RECT  3.255000  0.675000  3.425000 1.015000 ;
      RECT  3.255000  1.015000  3.460000 1.185000 ;
      RECT  3.290000  1.185000  3.460000 1.935000 ;
      RECT  3.290000  1.935000  5.075000 2.105000 ;
      RECT  3.460000  2.105000  3.630000 2.465000 ;
      RECT  3.680000  0.425000  3.850000 1.685000 ;
      RECT  4.300000  2.275000  4.630000 2.635000 ;
      RECT  4.445000  0.085000  4.775000 0.540000 ;
      RECT  4.565000  0.715000  5.145000 0.895000 ;
      RECT  4.565000  0.895000  4.735000 1.935000 ;
      RECT  4.905000  1.065000  5.075000 1.395000 ;
      RECT  4.905000  2.105000  5.075000 2.185000 ;
      RECT  4.905000  2.185000  5.275000 2.435000 ;
      RECT  4.975000  0.335000  5.315000 0.505000 ;
      RECT  4.975000  0.505000  5.145000 0.715000 ;
      RECT  5.245000  1.575000  5.495000 1.955000 ;
      RECT  5.325000  0.705000  5.975000 1.035000 ;
      RECT  5.325000  1.035000  5.495000 1.575000 ;
      RECT  5.470000  2.135000  5.835000 2.465000 ;
      RECT  5.485000  0.305000  6.335000 0.475000 ;
      RECT  5.665000  1.215000  7.375000 1.385000 ;
      RECT  5.665000  1.385000  5.835000 2.135000 ;
      RECT  6.005000  1.935000  7.165000 2.105000 ;
      RECT  6.005000  2.105000  6.175000 2.375000 ;
      RECT  6.165000  0.475000  6.335000 1.215000 ;
      RECT  6.285000  1.595000  7.715000 1.765000 ;
      RECT  6.410000  2.355000  6.740000 2.635000 ;
      RECT  6.915000  0.085000  7.245000 0.545000 ;
      RECT  6.995000  2.105000  7.165000 2.375000 ;
      RECT  7.205000  1.005000  7.375000 1.215000 ;
      RECT  7.375000  2.175000  7.745000 2.635000 ;
      RECT  7.455000  0.275000  7.785000 0.445000 ;
      RECT  7.455000  0.445000  7.715000 0.835000 ;
      RECT  7.455000  1.765000  7.715000 1.835000 ;
      RECT  7.455000  1.835000  8.140000 2.005000 ;
      RECT  7.545000  0.835000  7.715000 1.595000 ;
      RECT  7.885000  0.705000  8.095000 1.495000 ;
      RECT  7.885000  1.495000  8.520000 1.655000 ;
      RECT  7.885000  1.655000  8.870000 1.665000 ;
      RECT  7.970000  2.005000  8.140000 2.465000 ;
      RECT  8.005000  0.255000  8.915000 0.535000 ;
      RECT  8.310000  1.665000  8.870000 1.935000 ;
      RECT  8.310000  1.935000  8.840000 1.955000 ;
      RECT  8.320000  2.125000  9.190000 2.465000 ;
      RECT  8.405000  0.920000  8.575000 1.325000 ;
      RECT  8.745000  0.535000  8.915000 1.315000 ;
      RECT  8.745000  1.315000  9.210000 1.485000 ;
      RECT  9.015000  2.035000  9.210000 2.115000 ;
      RECT  9.015000  2.115000  9.190000 2.125000 ;
      RECT  9.040000  1.485000  9.210000 1.575000 ;
      RECT  9.040000  1.575000 10.205000 1.745000 ;
      RECT  9.040000  1.745000  9.210000 2.035000 ;
      RECT  9.085000  0.085000  9.255000 0.525000 ;
      RECT  9.125000  0.695000  9.655000 0.865000 ;
      RECT  9.125000  0.865000  9.295000 1.145000 ;
      RECT  9.360000  2.195000  9.610000 2.635000 ;
      RECT  9.485000  0.295000 10.515000 0.465000 ;
      RECT  9.485000  0.465000  9.655000 0.695000 ;
      RECT  9.780000  1.915000 10.545000 2.085000 ;
      RECT  9.780000  2.085000  9.950000 2.375000 ;
      RECT 10.120000  2.255000 10.450000 2.635000 ;
      RECT 10.345000  0.465000 10.515000 0.995000 ;
      RECT 10.345000  0.995000 11.020000 1.295000 ;
      RECT 10.375000  1.295000 11.020000 1.325000 ;
      RECT 10.375000  1.325000 10.545000 1.915000 ;
      RECT 10.720000  0.085000 10.890000 0.545000 ;
      RECT 10.720000  1.495000 10.970000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.675000  1.785000  0.845000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.145000  1.105000  1.315000 1.275000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.905000  1.105000  5.075000 1.275000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.325000  1.785000  5.495000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.405000  1.105000  8.575000 1.275000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.445000  1.785000  8.615000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
    LAYER met1 ;
      RECT 0.615000 1.755000 0.915000 1.800000 ;
      RECT 0.615000 1.800000 8.675000 1.940000 ;
      RECT 0.615000 1.940000 0.915000 1.985000 ;
      RECT 1.085000 1.075000 1.375000 1.120000 ;
      RECT 1.085000 1.120000 8.635000 1.260000 ;
      RECT 1.085000 1.260000 1.375000 1.305000 ;
      RECT 4.845000 1.075000 5.135000 1.120000 ;
      RECT 4.845000 1.260000 5.135000 1.305000 ;
      RECT 5.265000 1.755000 5.555000 1.800000 ;
      RECT 5.265000 1.940000 5.555000 1.985000 ;
      RECT 8.345000 1.075000 8.635000 1.120000 ;
      RECT 8.345000 1.260000 8.635000 1.305000 ;
      RECT 8.385000 1.755000 8.675000 1.800000 ;
      RECT 8.385000 1.940000 8.675000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfrtn_1
MACRO sky130_fd_sc_hd__nand3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.330000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.075000 2.160000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 1.075000 3.595000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 0.845000 1.445000 ;
        RECT 0.515000 1.445000 3.045000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 2.715000 1.665000 3.045000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.295000 2.105000 0.465000 ;
      RECT 0.090000  0.465000 0.345000 0.785000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.355000  0.635000 3.045000 0.905000 ;
      RECT 1.855000  1.835000 2.545000 2.635000 ;
      RECT 2.295000  0.085000 2.625000 0.465000 ;
      RECT 3.215000  0.085000 3.595000 0.885000 ;
      RECT 3.215000  1.445000 3.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__nand3_2
MACRO sky130_fd_sc_hd__nand3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 0.995000 1.755000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 0.765000 1.240000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.745000 0.330000 1.325000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.699000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 1.745000 0.595000 ;
        RECT 0.515000 0.595000 0.695000 1.495000 ;
        RECT 0.515000 1.495000 1.745000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.415000 0.595000 1.745000 0.825000 ;
        RECT 1.415000 1.665000 1.745000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.575000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 1.015000  1.835000 1.245000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__nand3_1
MACRO sky130_fd_sc_hd__nand3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.850000 1.075000 5.565000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.075000 3.540000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.700000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.445000 6.355000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 2.195000 1.665000 2.525000 2.465000 ;
        RECT 3.035000 1.665000 3.365000 2.465000 ;
        RECT 4.395000 0.655000 6.355000 0.905000 ;
        RECT 4.395000 1.665000 4.725000 2.465000 ;
        RECT 5.235000 1.665000 5.565000 2.465000 ;
        RECT 6.125000 0.905000 6.355000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 3.785000 0.905000 ;
      RECT 0.090000  1.445000 0.345000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.565000 ;
      RECT 0.935000  0.255000 1.265000 0.735000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.435000  0.085000 1.605000 0.565000 ;
      RECT 1.775000  0.655000 2.105000 0.735000 ;
      RECT 1.855000  1.835000 2.025000 2.635000 ;
      RECT 2.195000  0.255000 6.000000 0.485000 ;
      RECT 2.615000  0.655000 2.945000 0.735000 ;
      RECT 2.695000  1.835000 2.865000 2.635000 ;
      RECT 3.455000  0.655000 3.785000 0.735000 ;
      RECT 3.535000  1.835000 4.225000 2.635000 ;
      RECT 4.895000  1.835000 5.065000 2.635000 ;
      RECT 5.735000  1.835000 6.000000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__nand3_4
MACRO sky130_fd_sc_hd__dlygate4sd1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd1_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.555000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.410000 0.255000 2.700000 0.825000 ;
        RECT 2.440000 1.495000 2.700000 2.465000 ;
        RECT 2.530000 0.825000 2.700000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.785000 0.895000 2.005000 ;
      RECT 0.085000  2.005000 0.380000 2.465000 ;
      RECT 0.095000  0.255000 0.380000 0.715000 ;
      RECT 0.095000  0.715000 0.895000 0.885000 ;
      RECT 0.550000  0.085000 0.765000 0.545000 ;
      RECT 0.550000  2.175000 0.765000 2.635000 ;
      RECT 0.725000  0.885000 0.895000 0.995000 ;
      RECT 0.725000  0.995000 0.980000 1.325000 ;
      RECT 0.725000  1.325000 0.895000 1.785000 ;
      RECT 0.935000  0.255000 1.320000 0.545000 ;
      RECT 0.935000  2.175000 1.320000 2.465000 ;
      RECT 1.150000  0.545000 1.320000 1.075000 ;
      RECT 1.150000  1.075000 1.900000 1.275000 ;
      RECT 1.150000  1.275000 1.320000 2.175000 ;
      RECT 1.515000  0.255000 1.740000 0.735000 ;
      RECT 1.515000  0.735000 2.240000 0.905000 ;
      RECT 1.515000  1.575000 2.240000 1.745000 ;
      RECT 1.515000  1.745000 1.740000 2.430000 ;
      RECT 1.910000  0.085000 2.240000 0.565000 ;
      RECT 1.910000  1.915000 2.270000 2.635000 ;
      RECT 2.070000  0.905000 2.240000 0.995000 ;
      RECT 2.070000  0.995000 2.360000 1.325000 ;
      RECT 2.070000  1.325000 2.240000 1.575000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__dlygate4sd1_1
MACRO sky130_fd_sc_hd__a221oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.985000 1.075000 4.480000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.435000 1.075000 3.765000 1.445000 ;
        RECT 3.435000 1.445000 4.820000 1.615000 ;
        RECT 4.650000 1.075000 5.435000 1.275000 ;
        RECT 4.650000 1.275000 4.820000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.075000 2.765000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.075000 2.040000 1.445000 ;
        RECT 1.505000 1.445000 3.265000 1.615000 ;
        RECT 2.935000 1.075000 3.265000 1.445000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.420000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 0.305000 0.855000 0.725000 ;
        RECT 0.525000 0.725000 4.395000 0.865000 ;
        RECT 0.605000 0.865000 4.395000 0.905000 ;
        RECT 0.605000 0.905000 0.855000 2.125000 ;
        RECT 2.285000 0.645000 2.635000 0.725000 ;
        RECT 4.065000 0.645000 4.395000 0.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.090000  1.795000 0.435000 2.295000 ;
      RECT 0.090000  2.295000 1.275000 2.465000 ;
      RECT 0.105000  0.085000 0.355000 0.895000 ;
      RECT 1.025000  0.085000 1.715000 0.555000 ;
      RECT 1.025000  1.495000 1.275000 1.785000 ;
      RECT 1.025000  1.785000 3.015000 1.955000 ;
      RECT 1.025000  1.955000 1.275000 2.295000 ;
      RECT 1.505000  2.125000 1.755000 2.295000 ;
      RECT 1.505000  2.295000 3.475000 2.465000 ;
      RECT 1.885000  0.255000 3.055000 0.475000 ;
      RECT 1.925000  1.955000 2.175000 2.125000 ;
      RECT 2.345000  2.125000 2.595000 2.295000 ;
      RECT 2.765000  1.955000 3.015000 2.125000 ;
      RECT 3.225000  1.785000 5.195000 1.955000 ;
      RECT 3.225000  1.955000 3.475000 2.295000 ;
      RECT 3.270000  0.085000 3.440000 0.555000 ;
      RECT 3.645000  0.255000 4.815000 0.475000 ;
      RECT 3.685000  2.125000 3.935000 2.635000 ;
      RECT 4.105000  1.955000 4.355000 2.465000 ;
      RECT 4.525000  2.125000 4.775000 2.635000 ;
      RECT 4.565000  0.475000 4.815000 0.905000 ;
      RECT 4.985000  0.085000 5.155000 0.905000 ;
      RECT 4.990000  1.455000 5.195000 1.785000 ;
      RECT 4.990000  1.955000 5.195000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__a221oi_2
MACRO sky130_fd_sc_hd__a221oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 0.675000 2.200000 1.075000 ;
        RECT 1.945000 1.075000 2.275000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 0.995000 2.755000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 1.075000 1.695000 1.285000 ;
        RECT 1.415000 0.675000 1.695000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 1.075000 1.055000 1.285000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.435000 1.285000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.767000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.170000 0.255000 0.345000 0.735000 ;
        RECT 0.170000 0.735000 1.235000 0.905000 ;
        RECT 0.175000 1.455000 2.300000 1.495000 ;
        RECT 0.175000 1.495000 3.135000 1.625000 ;
        RECT 0.175000 1.625000 0.345000 2.465000 ;
        RECT 1.065000 0.255000 2.580000 0.505000 ;
        RECT 1.065000 0.505000 1.235000 0.735000 ;
        RECT 2.150000 1.625000 3.135000 1.665000 ;
        RECT 2.380000 0.505000 2.580000 0.655000 ;
        RECT 2.380000 0.655000 3.135000 0.825000 ;
        RECT 2.925000 0.825000 3.135000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.515000  0.085000 0.845000 0.565000 ;
      RECT 0.515000  1.795000 0.765000 2.295000 ;
      RECT 0.515000  2.295000 1.685000 2.465000 ;
      RECT 1.015000  1.795000 2.025000 1.835000 ;
      RECT 1.015000  1.835000 2.625000 2.045000 ;
      RECT 1.015000  2.045000 1.240000 2.125000 ;
      RECT 1.355000  2.255000 1.685000 2.295000 ;
      RECT 1.875000  2.215000 2.205000 2.635000 ;
      RECT 2.375000  2.045000 2.625000 2.465000 ;
      RECT 2.750000  0.085000 3.080000 0.485000 ;
      RECT 2.795000  1.875000 3.125000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a221oi_1
MACRO sky130_fd_sc_hd__a221oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.475000 1.075000 7.885000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.965000 1.075000 6.295000 1.445000 ;
        RECT 5.965000 1.445000 8.265000 1.615000 ;
        RECT 8.095000 1.075000 9.575000 1.275000 ;
        RECT 8.095000 1.275000 8.265000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.935000 0.995000 5.285000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.415000 0.995000 3.765000 1.325000 ;
        RECT 3.595000 1.325000 3.765000 1.445000 ;
        RECT 3.595000 1.445000 5.795000 1.615000 ;
        RECT 5.465000 1.075000 5.795000 1.445000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.335000 1.275000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 1.705000 0.905000 ;
        RECT 0.575000 1.445000 1.705000 1.615000 ;
        RECT 0.575000 1.615000 0.825000 2.125000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 1.415000 1.615000 1.665000 2.125000 ;
        RECT 1.505000 0.905000 1.705000 1.095000 ;
        RECT 1.505000 1.095000 3.245000 1.275000 ;
        RECT 1.505000 1.275000 1.705000 1.445000 ;
        RECT 3.075000 0.645000 5.680000 0.735000 ;
        RECT 3.075000 0.735000 7.765000 0.820000 ;
        RECT 3.075000 0.820000 3.245000 1.095000 ;
        RECT 5.510000 0.820000 6.460000 0.905000 ;
        RECT 6.290000 0.645000 7.765000 0.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.090000  1.445000 0.405000 2.295000 ;
      RECT 0.090000  2.295000 2.125000 2.465000 ;
      RECT 0.115000  0.085000 0.365000 0.895000 ;
      RECT 0.995000  1.785000 1.245000 2.295000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.875000  0.085000 2.045000 0.645000 ;
      RECT 1.875000  0.645000 2.905000 0.925000 ;
      RECT 1.875000  1.445000 3.030000 1.615000 ;
      RECT 1.875000  1.615000 2.125000 2.295000 ;
      RECT 2.235000  0.255000 5.585000 0.425000 ;
      RECT 2.235000  0.425000 2.610000 0.475000 ;
      RECT 2.315000  1.795000 2.565000 2.215000 ;
      RECT 2.315000  2.215000 6.005000 2.465000 ;
      RECT 2.735000  0.595000 2.905000 0.645000 ;
      RECT 2.735000  1.615000 3.030000 1.835000 ;
      RECT 2.735000  1.835000 5.585000 2.045000 ;
      RECT 3.035000  0.425000 5.585000 0.475000 ;
      RECT 5.755000  1.785000 8.605000 2.045000 ;
      RECT 5.755000  2.045000 6.005000 2.215000 ;
      RECT 5.835000  0.085000 6.005000 0.555000 ;
      RECT 6.175000  0.255000 8.185000 0.475000 ;
      RECT 6.175000  2.215000 8.185000 2.635000 ;
      RECT 7.935000  0.475000 8.185000 0.725000 ;
      RECT 7.935000  0.725000 9.025000 0.905000 ;
      RECT 8.355000  0.085000 8.525000 0.555000 ;
      RECT 8.355000  2.045000 8.525000 2.465000 ;
      RECT 8.435000  1.445000 9.405000 1.615000 ;
      RECT 8.435000  1.615000 8.605000 1.785000 ;
      RECT 8.695000  0.255000 9.025000 0.725000 ;
      RECT 8.775000  1.795000 8.945000 2.635000 ;
      RECT 9.155000  1.615000 9.405000 2.465000 ;
      RECT 9.195000  0.085000 9.365000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__a221oi_4
MACRO sky130_fd_sc_hd__fahcon_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fahcon_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.42000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 1.075000 1.340000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.937500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 0.710000 1.780000 1.325000 ;
      LAYER mcon ;
        RECT 1.525000 0.765000 1.695000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.265000 0.645000 4.515000 1.325000 ;
      LAYER mcon ;
        RECT 4.310000 0.765000 4.480000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465000 0.735000 1.755000 0.780000 ;
        RECT 1.465000 0.780000 4.540000 0.920000 ;
        RECT 1.465000 0.920000 1.755000 0.965000 ;
        RECT 4.250000 0.735000 4.540000 0.780000 ;
        RECT 4.250000 0.920000 4.540000 0.965000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.493500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.530000 1.075000 10.975000 1.275000 ;
    END
  END CI
  PIN COUT_N
    ANTENNADIFFAREA  0.402800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.610000 0.755000 6.935000 0.925000 ;
        RECT 6.610000 0.925000 6.880000 1.675000 ;
        RECT 6.710000 1.675000 6.880000 1.785000 ;
        RECT 6.765000 0.595000 6.935000 0.755000 ;
    END
  END COUT_N
  PIN SUM
    ANTENNADIFFAREA  0.463750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995000 0.255000 12.335000 0.825000 ;
        RECT 12.010000 1.785000 12.335000 2.465000 ;
        RECT 12.135000 0.825000 12.335000 1.785000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.610000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.085000  0.735000  0.430000 0.805000 ;
      RECT  0.085000  0.805000  0.255000 1.500000 ;
      RECT  0.085000  1.500000  0.440000 1.840000 ;
      RECT  0.085000  1.840000  1.110000 2.010000 ;
      RECT  0.085000  2.010000  0.430000 2.465000 ;
      RECT  0.100000  0.255000  0.430000 0.735000 ;
      RECT  0.425000  0.995000  0.780000 1.325000 ;
      RECT  0.600000  2.180000  0.770000 2.635000 ;
      RECT  0.610000  0.735000  1.325000 0.905000 ;
      RECT  0.610000  0.905000  0.780000 0.995000 ;
      RECT  0.610000  1.325000  0.780000 1.500000 ;
      RECT  0.610000  1.500000  1.450000 1.670000 ;
      RECT  0.630000  0.085000  0.800000 0.545000 ;
      RECT  0.940000  2.010000  1.110000 2.215000 ;
      RECT  0.940000  2.215000  2.545000 2.295000 ;
      RECT  0.940000  2.295000  3.540000 2.385000 ;
      RECT  0.995000  0.255000  3.410000 0.465000 ;
      RECT  0.995000  0.465000  1.325000 0.735000 ;
      RECT  1.280000  1.670000  1.450000 1.875000 ;
      RECT  1.280000  1.875000  2.920000 2.045000 ;
      RECT  1.965000  0.635000  2.470000 1.705000 ;
      RECT  2.375000  2.385000  3.540000 2.465000 ;
      RECT  2.640000  0.655000  3.025000 0.735000 ;
      RECT  2.640000  0.735000  3.160000 0.755000 ;
      RECT  2.640000  0.755000  3.750000 0.905000 ;
      RECT  2.640000  1.075000  2.975000 1.160000 ;
      RECT  2.640000  1.160000  3.100000 1.615000 ;
      RECT  3.055000  0.905000  3.750000 0.925000 ;
      RECT  3.240000  0.465000  3.410000 0.585000 ;
      RECT  3.270000  0.925000  3.440000 2.295000 ;
      RECT  3.580000  0.255000  4.595000 0.425000 ;
      RECT  3.580000  0.425000  3.750000 0.755000 ;
      RECT  3.725000  1.150000  4.095000 1.320000 ;
      RECT  3.725000  1.320000  3.895000 2.295000 ;
      RECT  3.725000  2.295000  5.100000 2.465000 ;
      RECT  3.925000  0.595000  4.095000 1.150000 ;
      RECT  4.210000  1.755000  4.380000 2.095000 ;
      RECT  4.265000  0.425000  4.595000 0.475000 ;
      RECT  4.700000  1.385000  5.180000 1.725000 ;
      RECT  4.840000  0.510000  5.030000 0.995000 ;
      RECT  4.840000  0.995000  5.180000 1.385000 ;
      RECT  4.875000  1.895000  6.005000 2.065000 ;
      RECT  4.875000  2.065000  5.100000 2.295000 ;
      RECT  5.200000  0.085000  5.530000 0.805000 ;
      RECT  5.270000  2.235000  5.600000 2.635000 ;
      RECT  5.645000  1.555000  6.380000 1.725000 ;
      RECT  5.700000  0.380000  5.980000 0.815000 ;
      RECT  5.810000  0.815000  5.980000 1.555000 ;
      RECT  5.835000  2.065000  6.005000 2.295000 ;
      RECT  5.835000  2.295000  7.960000 2.465000 ;
      RECT  6.150000  0.740000  6.435000 1.325000 ;
      RECT  6.210000  1.725000  6.380000 1.895000 ;
      RECT  6.210000  1.895000  6.540000 1.955000 ;
      RECT  6.210000  1.955000  7.220000 2.125000 ;
      RECT  6.265000  0.255000  7.700000 0.425000 ;
      RECT  6.265000  0.425000  6.595000 0.570000 ;
      RECT  7.050000  1.060000  7.280000 1.230000 ;
      RECT  7.050000  1.230000  7.220000 1.955000 ;
      RECT  7.110000  0.595000  7.360000 0.925000 ;
      RECT  7.110000  0.925000  7.280000 1.060000 ;
      RECT  7.390000  1.360000  7.620000 1.530000 ;
      RECT  7.390000  1.530000  7.560000 2.125000 ;
      RECT  7.450000  1.105000  7.700000 1.290000 ;
      RECT  7.450000  1.290000  7.620000 1.360000 ;
      RECT  7.530000  0.425000  7.700000 1.105000 ;
      RECT  7.790000  1.550000  8.045000 1.720000 ;
      RECT  7.790000  1.720000  7.960000 2.295000 ;
      RECT  7.875000  0.995000  8.045000 1.550000 ;
      RECT  7.935000  0.255000  9.450000 0.425000 ;
      RECT  7.935000  0.425000  8.270000 0.825000 ;
      RECT  8.230000  1.785000  8.400000 2.295000 ;
      RECT  8.230000  2.295000  9.950000 2.465000 ;
      RECT  8.440000  0.595000  8.900000 0.765000 ;
      RECT  8.440000  0.765000  8.610000 1.445000 ;
      RECT  8.440000  1.445000  8.740000 1.530000 ;
      RECT  8.440000  1.530000  8.900000 1.615000 ;
      RECT  8.570000  1.615000  8.900000 2.125000 ;
      RECT  8.780000  0.995000  9.110000 1.275000 ;
      RECT  9.070000  1.530000  9.450000 2.045000 ;
      RECT  9.070000  2.045000  9.420000 2.125000 ;
      RECT  9.280000  0.425000  9.450000 1.530000 ;
      RECT  9.620000  2.215000  9.950000 2.295000 ;
      RECT  9.650000  0.255000 10.020000 0.825000 ;
      RECT  9.650000  0.825000  9.820000 1.535000 ;
      RECT  9.650000  1.535000  9.950000 2.215000 ;
      RECT  9.990000  0.995000 10.360000 1.325000 ;
      RECT 10.120000  2.275000 10.455000 2.635000 ;
      RECT 10.190000  0.735000 10.920000 0.905000 ;
      RECT 10.190000  0.905000 10.360000 0.995000 ;
      RECT 10.190000  1.325000 10.360000 1.455000 ;
      RECT 10.190000  1.455000 10.835000 2.045000 ;
      RECT 10.200000  0.085000 10.370000 0.565000 ;
      RECT 10.540000  0.285000 10.920000 0.735000 ;
      RECT 10.625000  2.045000 10.835000 2.465000 ;
      RECT 11.085000  1.455000 11.415000 2.465000 ;
      RECT 11.165000  0.270000 11.335000 0.680000 ;
      RECT 11.165000  0.680000 11.415000 1.455000 ;
      RECT 11.535000  0.085000 11.825000 0.555000 ;
      RECT 11.585000  1.785000 11.840000 2.635000 ;
      RECT 11.655000  0.995000 11.965000 1.615000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.280000  1.785000  1.450000 1.955000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  1.105000  2.155000 1.275000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  2.930000  1.445000  3.100000 1.615000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.210000  1.785000  4.380000 1.955000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.770000  1.445000  4.940000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.150000  1.105000  6.320000 1.275000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.530000  0.765000  7.700000 0.935000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.450000  1.445000  8.620000 1.615000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.910000  1.105000  9.080000 1.275000 ;
      RECT  9.280000  1.785000  9.450000 1.955000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.190000  1.785000 10.360000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.230000  0.765000 11.400000 0.935000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 11.690000  1.445000 11.860000 1.615000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
    LAYER met1 ;
      RECT  1.195000 1.755000  1.510000 1.800000 ;
      RECT  1.195000 1.800000  4.440000 1.940000 ;
      RECT  1.195000 1.940000  1.510000 1.985000 ;
      RECT  1.925000 1.075000  2.215000 1.120000 ;
      RECT  1.925000 1.120000  9.140000 1.260000 ;
      RECT  1.925000 1.260000  2.215000 1.305000 ;
      RECT  2.845000 1.415000  3.160000 1.460000 ;
      RECT  2.845000 1.460000  5.000000 1.600000 ;
      RECT  2.845000 1.600000  3.160000 1.645000 ;
      RECT  4.150000 1.755000  4.440000 1.800000 ;
      RECT  4.150000 1.940000  4.440000 1.985000 ;
      RECT  4.710000 1.415000  5.000000 1.460000 ;
      RECT  4.710000 1.600000  5.000000 1.645000 ;
      RECT  6.090000 1.075000  6.380000 1.120000 ;
      RECT  6.090000 1.260000  6.380000 1.305000 ;
      RECT  7.470000 0.735000  7.760000 0.780000 ;
      RECT  7.470000 0.780000 11.460000 0.920000 ;
      RECT  7.470000 0.920000  7.760000 0.965000 ;
      RECT  8.390000 1.415000  8.680000 1.460000 ;
      RECT  8.390000 1.460000 11.920000 1.600000 ;
      RECT  8.390000 1.600000  8.680000 1.645000 ;
      RECT  8.850000 1.075000  9.140000 1.120000 ;
      RECT  8.850000 1.260000  9.140000 1.305000 ;
      RECT  9.195000 1.755000  9.510000 1.800000 ;
      RECT  9.195000 1.800000 10.420000 1.940000 ;
      RECT  9.195000 1.940000  9.510000 1.985000 ;
      RECT 10.130000 1.755000 10.420000 1.800000 ;
      RECT 10.130000 1.940000 10.420000 1.985000 ;
      RECT 11.170000 0.735000 11.460000 0.780000 ;
      RECT 11.170000 0.920000 11.460000 0.965000 ;
      RECT 11.630000 1.415000 11.920000 1.460000 ;
      RECT 11.630000 1.600000 11.920000 1.645000 ;
  END
END sky130_fd_sc_hd__fahcon_1
MACRO sky130_fd_sc_hd__o2111a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.830000 1.005000 4.515000 1.315000 ;
        RECT 4.310000 1.315000 4.515000 2.355000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.300000 0.995000 3.660000 1.325000 ;
        RECT 3.370000 1.325000 3.660000 2.370000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.680000 1.075000 3.100000 1.615000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 0.255000 2.390000 1.615000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.075000 1.835000 1.615000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.855000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.135000  0.085000 0.345000 0.885000 ;
      RECT 0.135000  1.495000 0.345000 2.635000 ;
      RECT 1.030000  0.715000 1.805000 0.885000 ;
      RECT 1.030000  0.885000 1.305000 1.785000 ;
      RECT 1.030000  1.785000 3.195000 2.025000 ;
      RECT 1.035000  0.085000 1.285000 0.545000 ;
      RECT 1.035000  2.195000 1.655000 2.635000 ;
      RECT 1.475000  0.255000 1.805000 0.715000 ;
      RECT 1.860000  2.025000 2.140000 2.465000 ;
      RECT 2.325000  2.255000 2.655000 2.635000 ;
      RECT 2.865000  0.255000 3.195000 0.625000 ;
      RECT 2.865000  0.625000 4.215000 0.825000 ;
      RECT 2.865000  2.025000 3.195000 2.465000 ;
      RECT 3.385000  0.085000 3.715000 0.455000 ;
      RECT 3.885000  0.255000 4.215000 0.625000 ;
      RECT 3.885000  1.495000 4.140000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__o2111a_2
MACRO sky130_fd_sc_hd__o2111a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.705000 1.075000 4.035000 1.660000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.050000 1.075000 3.535000 1.325000 ;
        RECT 3.350000 1.325000 3.535000 2.415000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.390000 2.690000 0.995000 ;
        RECT 2.445000 0.995000 2.705000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 0.390000 2.195000 1.325000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.265000 1.075000 1.745000 1.325000 ;
        RECT 1.535000 0.390000 1.745000 1.075000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.255000 0.355000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.525000  0.995000 0.865000 1.325000 ;
      RECT 0.525000  1.835000 1.335000 2.635000 ;
      RECT 0.535000  0.085000 0.845000 0.565000 ;
      RECT 0.695000  0.735000 1.365000 0.905000 ;
      RECT 0.695000  0.905000 0.865000 0.995000 ;
      RECT 0.695000  1.325000 0.865000 1.495000 ;
      RECT 0.695000  1.495000 3.180000 1.665000 ;
      RECT 1.025000  0.255000 1.365000 0.735000 ;
      RECT 1.505000  1.665000 1.835000 2.465000 ;
      RECT 2.020000  1.835000 2.760000 2.635000 ;
      RECT 2.870000  0.255000 3.160000 0.705000 ;
      RECT 2.870000  0.705000 4.055000 0.875000 ;
      RECT 2.930000  1.665000 3.180000 2.465000 ;
      RECT 3.330000  0.085000 3.620000 0.535000 ;
      RECT 3.730000  1.835000 4.055000 2.635000 ;
      RECT 3.790000  0.255000 4.055000 0.705000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o2111a_1
MACRO sky130_fd_sc_hd__o2111a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.890000 1.075000 4.485000 1.245000 ;
        RECT 4.130000 1.245000 4.485000 1.320000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.135000 1.075000 3.600000 1.245000 ;
        RECT 3.145000 1.245000 3.600000 1.320000 ;
        RECT 3.305000 1.320000 3.600000 1.490000 ;
        RECT 3.305000 1.490000 4.825000 1.660000 ;
        RECT 4.655000 1.075000 4.985000 1.320000 ;
        RECT 4.655000 1.320000 4.825000 1.490000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775000 1.075000 2.215000 1.320000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.150000 0.995000 1.395000 1.490000 ;
        RECT 1.150000 1.490000 2.660000 1.660000 ;
        RECT 2.445000 1.080000 2.820000 1.320000 ;
        RECT 2.445000 1.320000 2.660000 1.490000 ;
        RECT 2.490000 1.075000 2.820000 1.080000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.995000 0.340000 1.655000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.962500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.650000 0.255000 5.875000 0.695000 ;
        RECT 5.650000 0.695000 7.275000 0.865000 ;
        RECT 5.755000 1.495000 7.275000 1.665000 ;
        RECT 5.755000 1.665000 5.925000 2.465000 ;
        RECT 6.545000 0.255000 6.745000 0.695000 ;
        RECT 6.585000 1.665000 6.775000 2.465000 ;
        RECT 7.005000 0.865000 7.275000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.090000  1.835000 5.550000 2.000000 ;
      RECT 0.090000  2.000000 5.065000 2.005000 ;
      RECT 0.090000  2.005000 0.345000 2.465000 ;
      RECT 0.100000  0.255000 2.940000 0.485000 ;
      RECT 0.100000  0.485000 0.345000 0.825000 ;
      RECT 0.515000  0.655000 0.860000 1.830000 ;
      RECT 0.515000  1.830000 5.550000 1.835000 ;
      RECT 0.515000  2.175000 0.845000 2.635000 ;
      RECT 1.015000  2.005000 1.230000 2.465000 ;
      RECT 1.400000  2.175000 1.625000 2.635000 ;
      RECT 1.720000  0.655000 4.795000 0.885000 ;
      RECT 1.795000  2.005000 2.025000 2.465000 ;
      RECT 2.195000  2.175000 2.525000 2.635000 ;
      RECT 2.695000  2.005000 3.285000 2.465000 ;
      RECT 3.110000  0.085000 3.440000 0.485000 ;
      RECT 3.610000  0.255000 3.825000 0.655000 ;
      RECT 3.805000  2.180000 4.135000 2.635000 ;
      RECT 3.995000  0.085000 4.365000 0.485000 ;
      RECT 4.535000  0.255000 4.795000 0.655000 ;
      RECT 4.775000  2.005000 5.065000 2.465000 ;
      RECT 5.035000  0.085000 5.300000 0.545000 ;
      RECT 5.245000  2.170000 5.585000 2.635000 ;
      RECT 5.380000  1.075000 6.760000 1.320000 ;
      RECT 5.380000  1.320000 5.550000 1.830000 ;
      RECT 6.075000  0.085000 6.375000 0.525000 ;
      RECT 6.095000  1.835000 6.415000 2.635000 ;
      RECT 6.915000  0.085000 7.275000 0.525000 ;
      RECT 6.945000  1.835000 7.270000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__o2111a_4
MACRO sky130_fd_sc_hd__o311ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 1.105000 1.315000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275000 1.055000 2.155000 1.315000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 1.055000 3.075000 1.315000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.055000 4.385000 1.315000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.085000 1.055000 5.895000 1.315000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.551000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415000 1.485000 5.895000 1.725000 ;
        RECT 2.415000 1.725000 2.665000 2.125000 ;
        RECT 3.335000 1.725000 3.505000 2.465000 ;
        RECT 4.515000 1.725000 4.825000 2.465000 ;
        RECT 4.555000 0.655000 5.895000 0.885000 ;
        RECT 4.555000 0.885000 4.915000 1.485000 ;
        RECT 5.495000 1.725000 5.895000 2.465000 ;
        RECT 5.515000 0.255000 5.895000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.255000 0.485000 0.655000 ;
      RECT 0.085000  0.655000 4.385000 0.885000 ;
      RECT 0.085000  1.485000 2.225000 1.725000 ;
      RECT 0.085000  1.725000 0.465000 2.465000 ;
      RECT 0.635000  1.895000 0.965000 2.635000 ;
      RECT 0.655000  0.085000 0.985000 0.485000 ;
      RECT 1.135000  1.725000 1.305000 2.465000 ;
      RECT 1.155000  0.255000 1.325000 0.655000 ;
      RECT 1.475000  1.895000 1.805000 2.295000 ;
      RECT 1.475000  2.295000 3.165000 2.465000 ;
      RECT 1.495000  0.085000 1.825000 0.485000 ;
      RECT 1.975000  1.725000 2.225000 2.125000 ;
      RECT 1.995000  0.255000 2.165000 0.655000 ;
      RECT 2.335000  0.085000 3.105000 0.485000 ;
      RECT 2.835000  1.895000 3.165000 2.295000 ;
      RECT 3.275000  0.255000 3.445000 0.655000 ;
      RECT 3.615000  0.255000 5.345000 0.485000 ;
      RECT 3.675000  1.895000 4.345000 2.635000 ;
      RECT 4.995000  1.895000 5.325000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__o311ai_2
MACRO sky130_fd_sc_hd__o311ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.780000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.995000 1.260000 2.465000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.430000 0.995000 1.780000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.320000 2.200000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.830000 0.995000 3.135000 1.325000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.942000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.430000 1.495000 3.135000 1.665000 ;
        RECT 1.430000 1.665000 1.980000 2.465000 ;
        RECT 2.445000 0.255000 3.135000 0.825000 ;
        RECT 2.445000 0.825000 2.660000 1.495000 ;
        RECT 2.650000 1.665000 3.135000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.570000 0.825000 ;
      RECT 0.085000  1.495000 0.780000 2.635000 ;
      RECT 0.740000  0.255000 0.910000 0.655000 ;
      RECT 0.740000  0.655000 1.750000 0.825000 ;
      RECT 1.080000  0.085000 1.410000 0.485000 ;
      RECT 1.580000  0.255000 1.750000 0.655000 ;
      RECT 2.150000  1.835000 2.480000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o311ai_1
MACRO sky130_fd_sc_hd__o311ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 1.775000 1.315000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.055000 3.615000 1.315000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 1.055000 5.885000 1.315000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055000 1.055000 7.695000 1.315000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.865000 1.055000 9.090000 1.315000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.241000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.055000 1.485000 9.575000 1.725000 ;
        RECT 4.055000 1.725000 4.305000 2.115000 ;
        RECT 4.975000 1.725000 5.145000 2.115000 ;
        RECT 5.815000 1.725000 6.005000 2.465000 ;
        RECT 6.675000 1.725000 6.845000 2.465000 ;
        RECT 7.515000 1.725000 7.685000 2.465000 ;
        RECT 7.895000 0.655000 9.575000 0.885000 ;
        RECT 8.355000 1.725000 8.525000 2.465000 ;
        RECT 9.195000 1.725000 9.575000 2.465000 ;
        RECT 9.260000 0.885000 9.575000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125000 -0.085000 0.295000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.085000  0.085000 0.505000 0.885000 ;
      RECT 0.085000  1.485000 3.865000 1.725000 ;
      RECT 0.085000  1.725000 0.405000 2.465000 ;
      RECT 0.595000  1.895000 0.925000 2.635000 ;
      RECT 0.675000  0.255000 0.845000 0.655000 ;
      RECT 0.675000  0.655000 7.385000 0.885000 ;
      RECT 1.015000  0.085000 1.345000 0.485000 ;
      RECT 1.095000  1.725000 1.265000 2.465000 ;
      RECT 1.435000  1.895000 1.765000 2.635000 ;
      RECT 1.515000  0.255000 1.685000 0.655000 ;
      RECT 1.855000  0.085000 2.185000 0.485000 ;
      RECT 1.935000  1.725000 2.105000 2.465000 ;
      RECT 2.275000  1.895000 2.605000 2.295000 ;
      RECT 2.275000  2.295000 5.645000 2.465000 ;
      RECT 2.355000  0.255000 2.525000 0.655000 ;
      RECT 2.695000  0.085000 3.025000 0.485000 ;
      RECT 2.775000  1.725000 2.945000 2.115000 ;
      RECT 3.115000  1.895000 3.445000 2.295000 ;
      RECT 3.195000  0.255000 3.365000 0.655000 ;
      RECT 3.535000  0.085000 3.885000 0.485000 ;
      RECT 3.615000  1.725000 3.865000 2.115000 ;
      RECT 4.055000  0.255000 4.225000 0.655000 ;
      RECT 4.395000  0.085000 4.725000 0.485000 ;
      RECT 4.475000  1.895000 4.805000 2.295000 ;
      RECT 4.895000  0.255000 5.065000 0.655000 ;
      RECT 5.235000  0.085000 5.585000 0.485000 ;
      RECT 5.315000  1.895000 5.645000 2.295000 ;
      RECT 5.755000  0.255000 9.575000 0.485000 ;
      RECT 6.175000  1.895000 6.505000 2.635000 ;
      RECT 7.015000  1.895000 7.345000 2.635000 ;
      RECT 7.555000  0.485000 7.725000 0.885000 ;
      RECT 7.855000  1.895000 8.185000 2.635000 ;
      RECT 8.695000  1.895000 9.025000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__o311ai_4
MACRO sky130_fd_sc_hd__o311ai_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.570000 0.995000 ;
        RECT 0.085000 0.995000 0.780000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.995000 1.260000 2.465000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.430000 0.995000 1.780000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.260000 2.200000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.830000 0.765000 3.135000 1.325000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.604000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.430000 1.495000 3.135000 1.665000 ;
        RECT 1.430000 1.665000 1.980000 2.465000 ;
        RECT 2.445000 0.255000 3.135000 0.595000 ;
        RECT 2.445000 0.595000 2.660000 1.495000 ;
        RECT 2.650000 1.665000 3.135000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.570000 0.595000 ;
      RECT 0.085000  1.795000 0.780000 2.635000 ;
      RECT 0.740000  0.255000 0.910000 0.655000 ;
      RECT 0.740000  0.655000 1.750000 0.825000 ;
      RECT 1.080000  0.085000 1.410000 0.485000 ;
      RECT 1.580000  0.255000 1.750000 0.655000 ;
      RECT 2.150000  1.835000 2.480000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o311ai_0
MACRO sky130_fd_sc_hd__dlygate4sd2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.625000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.570000 0.255000 3.135000 0.825000 ;
        RECT 2.570000 1.495000 3.135000 2.465000 ;
        RECT 2.675000 0.825000 3.135000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.255000 0.485000 0.715000 ;
      RECT 0.085000  0.715000 1.030000 0.885000 ;
      RECT 0.085000  1.785000 1.030000 2.005000 ;
      RECT 0.085000  2.005000 0.485000 2.465000 ;
      RECT 0.655000  0.085000 0.925000 0.545000 ;
      RECT 0.655000  2.175000 0.925000 2.635000 ;
      RECT 0.795000  0.885000 1.030000 0.995000 ;
      RECT 0.795000  0.995000 1.085000 1.325000 ;
      RECT 0.795000  1.325000 1.030000 1.785000 ;
      RECT 1.155000  0.255000 1.425000 0.585000 ;
      RECT 1.155000  2.135000 1.425000 2.465000 ;
      RECT 1.255000  0.585000 1.425000 1.055000 ;
      RECT 1.255000  1.055000 2.030000 1.615000 ;
      RECT 1.255000  1.615000 1.425000 2.135000 ;
      RECT 1.615000  0.255000 1.875000 0.715000 ;
      RECT 1.615000  0.715000 2.400000 0.885000 ;
      RECT 1.615000  1.785000 2.400000 2.005000 ;
      RECT 1.615000  2.005000 1.875000 2.465000 ;
      RECT 2.075000  0.085000 2.400000 0.545000 ;
      RECT 2.075000  2.175000 2.400000 2.635000 ;
      RECT 2.200000  0.885000 2.400000 0.995000 ;
      RECT 2.200000  0.995000 2.505000 1.325000 ;
      RECT 2.200000  1.325000 2.400000 1.785000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__dlygate4sd2_1
MACRO sky130_fd_sc_hd__xor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.525000 1.075000 8.935000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705000 0.995000 7.875000 1.445000 ;
        RECT 7.705000 1.445000 8.285000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.880000 0.995000 3.515000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.350000 0.765000 0.660000 ;
        RECT 0.595000 0.660000 1.605000 0.830000 ;
        RECT 0.595000 0.830000 1.535000 0.925000 ;
        RECT 0.695000 1.440000 1.420000 1.455000 ;
        RECT 0.695000 1.455000 1.705000 2.045000 ;
        RECT 0.695000 2.045000 0.865000 2.465000 ;
        RECT 1.105000 0.925000 1.420000 1.440000 ;
        RECT 1.435000 0.350000 1.605000 0.660000 ;
        RECT 1.535000 2.045000 1.705000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 0.175000  0.085000  0.345000 0.545000 ;
        RECT 0.935000  0.085000  1.265000 0.465000 ;
        RECT 1.855000  0.085000  2.025000 0.525000 ;
        RECT 4.950000  0.085000  5.120000 0.885000 ;
        RECT 8.995000  0.085000  9.165000 0.565000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
        RECT 8.885000 -0.085000 9.055000 0.085000 ;
        RECT 9.345000 -0.085000 9.515000 0.085000 ;
        RECT 9.805000 -0.085000 9.975000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.235000 -0.085000 0.405000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 0.275000 2.135000  0.445000 2.635000 ;
        RECT 1.035000 2.215000  1.365000 2.635000 ;
        RECT 1.875000 2.215000  2.205000 2.635000 ;
        RECT 4.705000 2.235000  5.035000 2.635000 ;
        RECT 8.915000 2.275000  9.245000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
        RECT 8.885000 2.635000 9.055000 2.805000 ;
        RECT 9.345000 2.635000 9.515000 2.805000 ;
        RECT 9.805000 2.635000 9.975000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.820000 0.965000 2.045000 1.325000 ;
      RECT 1.875000 0.695000 2.365000 0.865000 ;
      RECT 1.875000 0.865000 2.045000 0.965000 ;
      RECT 1.875000 1.325000 2.045000 1.875000 ;
      RECT 1.875000 1.875000 2.545000 2.045000 ;
      RECT 2.195000 0.255000 3.760000 0.425000 ;
      RECT 2.195000 0.425000 2.365000 0.695000 ;
      RECT 2.370000 1.535000 3.855000 1.705000 ;
      RECT 2.375000 2.045000 2.545000 2.235000 ;
      RECT 2.375000 2.235000 3.915000 2.405000 ;
      RECT 2.540000 0.595000 2.710000 1.535000 ;
      RECT 2.890000 1.895000 4.195000 2.065000 ;
      RECT 2.990000 0.655000 4.100000 0.825000 ;
      RECT 3.410000 0.425000 3.760000 0.455000 ;
      RECT 3.685000 0.995000 4.055000 1.325000 ;
      RECT 3.685000 1.325000 3.855000 1.535000 ;
      RECT 3.930000 0.255000 4.780000 0.425000 ;
      RECT 3.930000 0.425000 4.100000 0.655000 ;
      RECT 4.025000 1.525000 4.555000 1.695000 ;
      RECT 4.025000 1.695000 4.195000 1.895000 ;
      RECT 4.130000 2.235000 4.535000 2.405000 ;
      RECT 4.270000 0.595000 4.440000 1.375000 ;
      RECT 4.270000 1.375000 4.555000 1.525000 ;
      RECT 4.365000 1.895000 5.540000 2.065000 ;
      RECT 4.365000 2.065000 4.535000 2.235000 ;
      RECT 4.610000 0.425000 4.780000 1.035000 ;
      RECT 4.610000 1.035000 4.865000 1.040000 ;
      RECT 4.610000 1.040000 4.880000 1.045000 ;
      RECT 4.610000 1.045000 4.890000 1.050000 ;
      RECT 4.610000 1.050000 4.895000 1.205000 ;
      RECT 4.725000 1.205000 4.895000 1.895000 ;
      RECT 5.125000 1.445000 5.540000 1.715000 ;
      RECT 5.300000 0.415000 5.540000 1.445000 ;
      RECT 5.370000 2.065000 5.540000 2.275000 ;
      RECT 5.370000 2.275000 8.465000 2.445000 ;
      RECT 5.715000 0.265000 6.130000 0.485000 ;
      RECT 5.715000 0.485000 5.935000 0.595000 ;
      RECT 5.715000 0.595000 5.885000 2.105000 ;
      RECT 6.075000 0.720000 6.470000 0.825000 ;
      RECT 6.075000 0.825000 6.275000 0.890000 ;
      RECT 6.075000 0.890000 6.245000 2.275000 ;
      RECT 6.105000 0.655000 6.470000 0.720000 ;
      RECT 6.300000 0.320000 6.470000 0.655000 ;
      RECT 6.415000 1.445000 7.195000 1.615000 ;
      RECT 6.415000 1.615000 6.830000 2.045000 ;
      RECT 6.430000 0.995000 6.855000 1.270000 ;
      RECT 6.640000 0.630000 6.855000 0.995000 ;
      RECT 7.025000 0.255000 8.170000 0.425000 ;
      RECT 7.025000 0.425000 7.195000 1.445000 ;
      RECT 7.365000 0.595000 7.535000 1.935000 ;
      RECT 7.365000 1.935000 9.675000 2.105000 ;
      RECT 7.705000 0.425000 8.170000 0.465000 ;
      RECT 8.045000 0.730000 8.250000 0.945000 ;
      RECT 8.045000 0.945000 8.355000 1.275000 ;
      RECT 8.455000 1.495000 9.275000 1.705000 ;
      RECT 8.495000 0.295000 8.785000 0.735000 ;
      RECT 8.495000 0.735000 9.275000 0.750000 ;
      RECT 8.535000 0.750000 9.275000 0.905000 ;
      RECT 9.105000 0.905000 9.275000 0.995000 ;
      RECT 9.105000 0.995000 9.335000 1.325000 ;
      RECT 9.105000 1.325000 9.275000 1.495000 ;
      RECT 9.190000 1.875000 9.675000 1.935000 ;
      RECT 9.415000 0.255000 9.675000 0.585000 ;
      RECT 9.415000 2.105000 9.675000 2.465000 ;
      RECT 9.505000 0.585000 9.675000 1.875000 ;
    LAYER mcon ;
      RECT 4.385000 1.445000 4.555000 1.615000 ;
      RECT 5.305000 0.765000 5.475000 0.935000 ;
      RECT 5.765000 0.425000 5.935000 0.595000 ;
      RECT 6.685000 0.765000 6.855000 0.935000 ;
      RECT 6.685000 1.445000 6.855000 1.615000 ;
      RECT 8.065000 0.765000 8.235000 0.935000 ;
      RECT 8.525000 0.425000 8.695000 0.595000 ;
    LAYER met1 ;
      RECT 4.325000 1.415000 4.615000 1.460000 ;
      RECT 4.325000 1.460000 6.915000 1.600000 ;
      RECT 4.325000 1.600000 4.615000 1.645000 ;
      RECT 5.245000 0.735000 5.535000 0.780000 ;
      RECT 5.245000 0.780000 8.295000 0.920000 ;
      RECT 5.245000 0.920000 5.535000 0.965000 ;
      RECT 5.705000 0.395000 5.995000 0.440000 ;
      RECT 5.705000 0.440000 8.755000 0.580000 ;
      RECT 5.705000 0.580000 5.995000 0.625000 ;
      RECT 6.625000 0.735000 6.915000 0.780000 ;
      RECT 6.625000 0.920000 6.915000 0.965000 ;
      RECT 6.625000 1.415000 6.915000 1.460000 ;
      RECT 6.625000 1.600000 6.915000 1.645000 ;
      RECT 8.005000 0.735000 8.295000 0.780000 ;
      RECT 8.005000 0.920000 8.295000 0.965000 ;
      RECT 8.465000 0.395000 8.755000 0.440000 ;
      RECT 8.465000 0.580000 8.755000 0.625000 ;
  END
END sky130_fd_sc_hd__xor3_4
MACRO sky130_fd_sc_hd__xor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.965000 1.075000 8.375000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.145000 0.995000 7.315000 1.445000 ;
        RECT 7.145000 1.445000 7.725000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.320000 0.995000 2.955000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.660000 1.050000 0.925000 ;
        RECT 0.545000 0.925000 0.860000 1.440000 ;
        RECT 0.545000 1.440000 1.070000 2.045000 ;
        RECT 0.800000 0.350000 1.050000 0.660000 ;
        RECT 0.820000 2.045000 1.070000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.300000  0.085000 0.630000 0.465000 ;
      RECT 0.300000  2.215000 0.650000 2.635000 ;
      RECT 1.210000  0.995000 1.410000 1.325000 ;
      RECT 1.220000  0.085000 1.470000 0.525000 ;
      RECT 1.240000  0.695000 1.810000 0.865000 ;
      RECT 1.240000  0.865000 1.410000 0.995000 ;
      RECT 1.240000  1.325000 1.410000 1.875000 ;
      RECT 1.240000  1.875000 1.930000 2.045000 ;
      RECT 1.240000  2.215000 1.575000 2.635000 ;
      RECT 1.640000  0.255000 3.200000 0.425000 ;
      RECT 1.640000  0.425000 1.810000 0.695000 ;
      RECT 1.645000  1.535000 3.295000 1.705000 ;
      RECT 1.760000  2.045000 1.930000 2.235000 ;
      RECT 1.760000  2.235000 3.355000 2.405000 ;
      RECT 1.980000  0.595000 2.150000 1.535000 ;
      RECT 2.330000  1.895000 3.635000 2.065000 ;
      RECT 2.430000  0.655000 3.540000 0.825000 ;
      RECT 2.850000  0.425000 3.200000 0.455000 ;
      RECT 3.125000  0.995000 3.400000 1.325000 ;
      RECT 3.125000  1.325000 3.295000 1.535000 ;
      RECT 3.370000  0.255000 4.220000 0.425000 ;
      RECT 3.370000  0.425000 3.540000 0.655000 ;
      RECT 3.465000  1.525000 3.995000 1.695000 ;
      RECT 3.465000  1.695000 3.635000 1.895000 ;
      RECT 3.570000  2.235000 3.975000 2.405000 ;
      RECT 3.710000  0.595000 3.880000 1.375000 ;
      RECT 3.710000  1.375000 3.995000 1.525000 ;
      RECT 3.805000  1.895000 4.980000 2.065000 ;
      RECT 3.805000  2.065000 3.975000 2.235000 ;
      RECT 4.050000  0.425000 4.220000 1.035000 ;
      RECT 4.050000  1.035000 4.335000 1.205000 ;
      RECT 4.145000  2.235000 4.475000 2.635000 ;
      RECT 4.165000  1.205000 4.335000 1.895000 ;
      RECT 4.390000  0.085000 4.560000 0.865000 ;
      RECT 4.565000  1.445000 4.980000 1.715000 ;
      RECT 4.740000  0.415000 4.980000 1.445000 ;
      RECT 4.810000  2.065000 4.980000 2.275000 ;
      RECT 4.810000  2.275000 7.905000 2.445000 ;
      RECT 5.155000  0.265000 5.570000 0.485000 ;
      RECT 5.155000  0.485000 5.375000 0.595000 ;
      RECT 5.155000  0.595000 5.325000 2.105000 ;
      RECT 5.495000  0.720000 5.910000 0.825000 ;
      RECT 5.495000  0.825000 5.715000 0.890000 ;
      RECT 5.495000  0.890000 5.665000 2.275000 ;
      RECT 5.545000  0.655000 5.910000 0.720000 ;
      RECT 5.740000  0.320000 5.910000 0.655000 ;
      RECT 5.855000  1.445000 6.635000 1.615000 ;
      RECT 5.855000  1.615000 6.270000 2.045000 ;
      RECT 5.870000  0.995000 6.295000 1.270000 ;
      RECT 6.080000  0.630000 6.295000 0.995000 ;
      RECT 6.465000  0.255000 7.610000 0.425000 ;
      RECT 6.465000  0.425000 6.635000 1.445000 ;
      RECT 6.805000  0.595000 6.975000 1.935000 ;
      RECT 6.805000  1.935000 9.115000 2.105000 ;
      RECT 7.145000  0.425000 7.610000 0.465000 ;
      RECT 7.485000  0.730000 7.690000 0.945000 ;
      RECT 7.485000  0.945000 7.795000 1.275000 ;
      RECT 7.895000  1.495000 8.715000 1.705000 ;
      RECT 7.935000  0.295000 8.225000 0.735000 ;
      RECT 7.935000  0.735000 8.715000 0.750000 ;
      RECT 7.975000  0.750000 8.715000 0.905000 ;
      RECT 8.315000  2.275000 8.650000 2.635000 ;
      RECT 8.395000  0.085000 8.565000 0.565000 ;
      RECT 8.545000  0.905000 8.715000 0.995000 ;
      RECT 8.545000  0.995000 8.775000 1.325000 ;
      RECT 8.545000  1.325000 8.715000 1.495000 ;
      RECT 8.630000  1.875000 9.115000 1.935000 ;
      RECT 8.815000  0.255000 9.115000 0.585000 ;
      RECT 8.820000  2.105000 9.115000 2.465000 ;
      RECT 8.945000  0.585000 9.115000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  1.445000 3.995000 1.615000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  0.765000 4.915000 0.935000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  0.425000 5.375000 0.595000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  0.765000 6.295000 0.935000 ;
      RECT 6.125000  1.445000 6.295000 1.615000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  0.765000 7.675000 0.935000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  0.425000 8.135000 0.595000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 3.765000 1.415000 4.055000 1.460000 ;
      RECT 3.765000 1.460000 6.355000 1.600000 ;
      RECT 3.765000 1.600000 4.055000 1.645000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.780000 7.735000 0.920000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.145000 0.395000 5.435000 0.440000 ;
      RECT 5.145000 0.440000 8.195000 0.580000 ;
      RECT 5.145000 0.580000 5.435000 0.625000 ;
      RECT 6.065000 0.735000 6.355000 0.780000 ;
      RECT 6.065000 0.920000 6.355000 0.965000 ;
      RECT 6.065000 1.415000 6.355000 1.460000 ;
      RECT 6.065000 1.600000 6.355000 1.645000 ;
      RECT 7.445000 0.735000 7.735000 0.780000 ;
      RECT 7.445000 0.920000 7.735000 0.965000 ;
      RECT 7.905000 0.395000 8.195000 0.440000 ;
      RECT 7.905000 0.580000 8.195000 0.625000 ;
  END
END sky130_fd_sc_hd__xor3_2
MACRO sky130_fd_sc_hd__xor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.505000 1.075000 7.915000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.685000 0.995000 6.855000 1.445000 ;
        RECT 6.685000 1.445000 7.265000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.860000 0.995000 2.495000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.590000 0.925000 ;
        RECT 0.085000 0.925000 0.400000 1.440000 ;
        RECT 0.085000 1.440000 0.610000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.750000  0.995000 0.950000 1.325000 ;
      RECT 0.760000  0.085000 1.010000 0.525000 ;
      RECT 0.780000  0.695000 1.350000 0.865000 ;
      RECT 0.780000  0.865000 0.950000 0.995000 ;
      RECT 0.780000  1.325000 0.950000 1.875000 ;
      RECT 0.780000  1.875000 1.470000 2.045000 ;
      RECT 0.780000  2.215000 1.115000 2.635000 ;
      RECT 1.180000  0.255000 2.740000 0.425000 ;
      RECT 1.180000  0.425000 1.350000 0.695000 ;
      RECT 1.185000  1.535000 2.835000 1.705000 ;
      RECT 1.300000  2.045000 1.470000 2.235000 ;
      RECT 1.300000  2.235000 2.895000 2.405000 ;
      RECT 1.520000  0.595000 1.690000 1.535000 ;
      RECT 1.870000  1.895000 3.175000 2.065000 ;
      RECT 1.970000  0.655000 3.080000 0.825000 ;
      RECT 2.390000  0.425000 2.740000 0.455000 ;
      RECT 2.665000  0.995000 2.940000 1.325000 ;
      RECT 2.665000  1.325000 2.835000 1.535000 ;
      RECT 2.910000  0.255000 3.760000 0.425000 ;
      RECT 2.910000  0.425000 3.080000 0.655000 ;
      RECT 3.005000  1.525000 3.535000 1.695000 ;
      RECT 3.005000  1.695000 3.175000 1.895000 ;
      RECT 3.110000  2.235000 3.515000 2.405000 ;
      RECT 3.250000  0.595000 3.420000 1.375000 ;
      RECT 3.250000  1.375000 3.535000 1.525000 ;
      RECT 3.345000  1.895000 4.520000 2.065000 ;
      RECT 3.345000  2.065000 3.515000 2.235000 ;
      RECT 3.590000  0.425000 3.760000 1.035000 ;
      RECT 3.590000  1.035000 3.875000 1.205000 ;
      RECT 3.685000  2.235000 4.015000 2.635000 ;
      RECT 3.705000  1.205000 3.875000 1.895000 ;
      RECT 3.930000  0.085000 4.100000 0.865000 ;
      RECT 4.105000  1.445000 4.520000 1.715000 ;
      RECT 4.280000  0.415000 4.520000 1.445000 ;
      RECT 4.350000  2.065000 4.520000 2.275000 ;
      RECT 4.350000  2.275000 7.445000 2.445000 ;
      RECT 4.695000  0.265000 5.110000 0.485000 ;
      RECT 4.695000  0.485000 4.915000 0.595000 ;
      RECT 4.695000  0.595000 4.865000 2.105000 ;
      RECT 5.035000  0.720000 5.450000 0.825000 ;
      RECT 5.035000  0.825000 5.255000 0.890000 ;
      RECT 5.035000  0.890000 5.205000 2.275000 ;
      RECT 5.085000  0.655000 5.450000 0.720000 ;
      RECT 5.280000  0.320000 5.450000 0.655000 ;
      RECT 5.395000  1.445000 6.175000 1.615000 ;
      RECT 5.395000  1.615000 5.810000 2.045000 ;
      RECT 5.410000  0.995000 5.835000 1.270000 ;
      RECT 5.620000  0.630000 5.835000 0.995000 ;
      RECT 6.005000  0.255000 7.150000 0.425000 ;
      RECT 6.005000  0.425000 6.175000 1.445000 ;
      RECT 6.345000  0.595000 6.515000 1.935000 ;
      RECT 6.345000  1.935000 8.655000 2.105000 ;
      RECT 6.685000  0.425000 7.150000 0.465000 ;
      RECT 7.025000  0.730000 7.230000 0.945000 ;
      RECT 7.025000  0.945000 7.335000 1.275000 ;
      RECT 7.435000  1.495000 8.255000 1.705000 ;
      RECT 7.475000  0.295000 7.765000 0.735000 ;
      RECT 7.475000  0.735000 8.255000 0.750000 ;
      RECT 7.515000  0.750000 8.255000 0.905000 ;
      RECT 7.855000  2.275000 8.190000 2.635000 ;
      RECT 7.935000  0.085000 8.105000 0.565000 ;
      RECT 8.085000  0.905000 8.255000 0.995000 ;
      RECT 8.085000  0.995000 8.315000 1.325000 ;
      RECT 8.085000  1.325000 8.255000 1.495000 ;
      RECT 8.170000  1.875000 8.655000 1.935000 ;
      RECT 8.355000  0.255000 8.655000 0.585000 ;
      RECT 8.360000  2.105000 8.655000 2.465000 ;
      RECT 8.485000  0.585000 8.655000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  1.445000 3.535000 1.615000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  0.765000 4.455000 0.935000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  0.425000 4.915000 0.595000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  0.765000 5.835000 0.935000 ;
      RECT 5.665000  1.445000 5.835000 1.615000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  0.765000 7.215000 0.935000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  0.425000 7.675000 0.595000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
    LAYER met1 ;
      RECT 3.305000 1.415000 3.595000 1.460000 ;
      RECT 3.305000 1.460000 5.895000 1.600000 ;
      RECT 3.305000 1.600000 3.595000 1.645000 ;
      RECT 4.225000 0.735000 4.515000 0.780000 ;
      RECT 4.225000 0.780000 7.275000 0.920000 ;
      RECT 4.225000 0.920000 4.515000 0.965000 ;
      RECT 4.685000 0.395000 4.975000 0.440000 ;
      RECT 4.685000 0.440000 7.735000 0.580000 ;
      RECT 4.685000 0.580000 4.975000 0.625000 ;
      RECT 5.605000 0.735000 5.895000 0.780000 ;
      RECT 5.605000 0.920000 5.895000 0.965000 ;
      RECT 5.605000 1.415000 5.895000 1.460000 ;
      RECT 5.605000 1.600000 5.895000 1.645000 ;
      RECT 6.985000 0.735000 7.275000 0.780000 ;
      RECT 6.985000 0.920000 7.275000 0.965000 ;
      RECT 7.445000 0.395000 7.735000 0.440000 ;
      RECT 7.445000 0.580000 7.735000 0.625000 ;
  END
END sky130_fd_sc_hd__xor3_1
MACRO sky130_fd_sc_hd__maj3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__maj3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 0.995000 1.695000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.865000 0.995000 2.155000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.495000 ;
        RECT 0.425000 1.495000 3.070000 1.665000 ;
        RECT 2.415000 1.415000 3.070000 1.495000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.285000 0.255000 3.615000 0.905000 ;
        RECT 3.285000 1.495000 3.615000 2.465000 ;
        RECT 3.445000 0.905000 3.615000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.280000 0.525000 0.655000 ;
      RECT 0.085000  0.655000 3.105000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.835000 ;
      RECT 0.085000  1.835000 2.085000 2.005000 ;
      RECT 0.085000  2.005000 0.615000 2.465000 ;
      RECT 0.975000  0.085000 1.305000 0.485000 ;
      RECT 0.975000  2.175000 1.305000 2.635000 ;
      RECT 1.755000  0.255000 2.085000 0.655000 ;
      RECT 1.755000  2.005000 2.085000 2.465000 ;
      RECT 2.535000  1.835000 2.860000 2.635000 ;
      RECT 2.635000  0.085000 2.965000 0.485000 ;
      RECT 2.925000  0.825000 3.105000 1.075000 ;
      RECT 2.925000  1.075000 3.275000 1.245000 ;
      RECT 3.785000  0.085000 4.055000 0.905000 ;
      RECT 3.785000  1.495000 4.055000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__maj3_2
MACRO sky130_fd_sc_hd__maj3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__maj3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 0.995000 1.125000 1.325000 ;
        RECT 0.610000 1.325000 0.780000 2.460000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 0.995000 1.905000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415000 0.765000 2.755000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.602250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.255000 0.255000 3.595000 0.825000 ;
        RECT 3.255000 2.160000 3.595000 2.465000 ;
        RECT 3.265000 1.495000 3.595000 2.160000 ;
        RECT 3.370000 0.825000 3.595000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.135000  0.255000 0.395000 0.655000 ;
      RECT 0.135000  0.655000 2.245000 0.825000 ;
      RECT 0.135000  0.825000 0.395000 2.125000 ;
      RECT 0.875000  0.085000 1.205000 0.485000 ;
      RECT 0.955000  1.715000 1.205000 2.635000 ;
      RECT 1.655000  0.255000 1.985000 0.640000 ;
      RECT 1.655000  0.640000 2.245000 0.655000 ;
      RECT 1.655000  1.815000 2.245000 2.080000 ;
      RECT 2.075000  0.825000 2.245000 1.495000 ;
      RECT 2.075000  1.495000 3.095000 1.665000 ;
      RECT 2.075000  1.665000 2.245000 1.815000 ;
      RECT 2.545000  0.085000 2.880000 0.470000 ;
      RECT 2.555000  1.845000 2.885000 2.635000 ;
      RECT 2.925000  0.995000 3.200000 1.325000 ;
      RECT 2.925000  1.325000 3.095000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__maj3_1
MACRO sky130_fd_sc_hd__maj3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__maj3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.075000 1.450000 1.635000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 1.075000 2.290000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 0.890000 1.285000 ;
        RECT 0.720000 1.285000 0.890000 1.915000 ;
        RECT 0.720000 1.915000 1.790000 2.085000 ;
        RECT 1.620000 2.085000 1.790000 2.225000 ;
        RECT 1.620000 2.225000 2.630000 2.395000 ;
        RECT 2.460000 1.075000 2.945000 1.245000 ;
        RECT 2.460000 1.245000 2.630000 2.225000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375000 0.255000 3.705000 0.490000 ;
        RECT 3.375000 1.455000 4.975000 1.625000 ;
        RECT 3.375000 1.625000 3.705000 2.465000 ;
        RECT 3.455000 0.490000 3.705000 0.715000 ;
        RECT 3.455000 0.715000 4.975000 0.905000 ;
        RECT 4.215000 0.255000 4.545000 0.715000 ;
        RECT 4.215000 1.625000 4.545000 2.465000 ;
        RECT 4.715000 0.905000 4.975000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.255000 0.635000 0.660000 ;
      RECT 0.085000  0.660000 2.290000 0.715000 ;
      RECT 0.085000  0.715000 3.285000 0.885000 ;
      RECT 0.085000  0.885000 0.255000 1.455000 ;
      RECT 0.085000  1.455000 0.465000 2.465000 ;
      RECT 1.120000  0.085000 1.450000 0.490000 ;
      RECT 1.120000  2.255000 1.450000 2.635000 ;
      RECT 1.620000  0.885000 1.790000 1.545000 ;
      RECT 1.620000  1.545000 2.290000 1.745000 ;
      RECT 1.960000  0.255000 2.290000 0.660000 ;
      RECT 1.960000  1.745000 2.290000 2.055000 ;
      RECT 2.845000  1.455000 3.175000 2.635000 ;
      RECT 2.860000  0.085000 3.205000 0.545000 ;
      RECT 3.115000  0.885000 3.285000 1.075000 ;
      RECT 3.115000  1.075000 4.545000 1.285000 ;
      RECT 3.875000  0.085000 4.045000 0.545000 ;
      RECT 3.875000  1.795000 4.045000 2.635000 ;
      RECT 4.715000  0.085000 4.885000 0.545000 ;
      RECT 4.715000  1.795000 4.925000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__maj3_4
MACRO sky130_fd_sc_hd__sedfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.18000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.935000 0.255000 14.265000 2.420000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.700000 1.065000 12.145000 1.300000 ;
        RECT 11.700000 1.300000 12.030000 2.465000 ;
        RECT 11.815000 0.255000 12.145000 1.065000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 1.105000 6.215000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.105000 5.250000 1.615000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.180000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  4.885000 1.435000 ;
        RECT -0.190000 1.435000 15.370000 2.910000 ;
        RECT  7.200000 1.305000 15.370000 1.435000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 15.180000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.180000 0.085000 ;
      RECT  0.000000  2.635000 15.180000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.595000  0.255000  4.795000 0.645000 ;
      RECT  4.595000  0.645000  4.855000 0.825000 ;
      RECT  4.635000  2.210000  4.965000 2.465000 ;
      RECT  4.685000  0.825000  4.855000 1.785000 ;
      RECT  4.685000  1.785000  4.965000 2.210000 ;
      RECT  4.965000  0.255000  5.590000 0.515000 ;
      RECT  5.155000  1.835000  6.585000 2.005000 ;
      RECT  5.155000  2.005000  5.495000 2.465000 ;
      RECT  5.260000  0.515000  5.590000 0.935000 ;
      RECT  5.420000  0.935000  5.590000 1.835000 ;
      RECT  5.665000  2.175000  6.010000 2.635000 ;
      RECT  5.760000  0.085000  6.010000 0.905000 ;
      RECT  6.385000  1.355000  6.585000 1.835000 ;
      RECT  6.515000  0.255000  7.135000 0.565000 ;
      RECT  6.515000  0.565000  6.925000 1.185000 ;
      RECT  6.675000  2.150000  7.005000 2.465000 ;
      RECT  6.755000  1.185000  6.925000 1.865000 ;
      RECT  6.755000  1.865000  7.005000 2.150000 ;
      RECT  7.095000  1.125000  7.280000 1.720000 ;
      RECT  7.115000  0.735000  7.620000 0.955000 ;
      RECT  7.215000  2.175000  8.255000 2.375000 ;
      RECT  7.305000  0.255000  7.980000 0.565000 ;
      RECT  7.450000  0.955000  7.620000 1.655000 ;
      RECT  7.450000  1.655000  7.915000 2.005000 ;
      RECT  7.810000  0.565000  7.980000 1.315000 ;
      RECT  7.810000  1.315000  8.660000 1.485000 ;
      RECT  8.085000  1.485000  8.660000 1.575000 ;
      RECT  8.085000  1.575000  8.255000 2.175000 ;
      RECT  8.170000  0.765000  9.235000 1.045000 ;
      RECT  8.170000  1.045000  9.745000 1.065000 ;
      RECT  8.170000  1.065000  8.370000 1.095000 ;
      RECT  8.245000  0.085000  8.640000 0.560000 ;
      RECT  8.425000  1.835000  8.660000 2.635000 ;
      RECT  8.490000  1.245000  8.660000 1.315000 ;
      RECT  8.830000  0.255000  9.235000 0.765000 ;
      RECT  8.830000  1.065000  9.745000 1.375000 ;
      RECT  8.830000  1.375000  9.160000 2.465000 ;
      RECT  9.370000  2.105000  9.660000 2.635000 ;
      RECT  9.465000  0.085000  9.740000 0.615000 ;
      RECT 10.090000  1.245000 10.280000 1.965000 ;
      RECT 10.225000  2.165000 11.190000 2.355000 ;
      RECT 10.305000  0.705000 10.770000 1.035000 ;
      RECT 10.325000  0.330000 11.190000 0.535000 ;
      RECT 10.450000  1.035000 10.770000 1.995000 ;
      RECT 10.940000  0.535000 11.190000 2.165000 ;
      RECT 11.360000  1.495000 11.530000 2.635000 ;
      RECT 11.395000  0.085000 11.645000 0.900000 ;
      RECT 12.200000  1.465000 12.450000 2.635000 ;
      RECT 12.315000  0.085000 12.565000 0.900000 ;
      RECT 12.620000  1.575000 12.850000 2.010000 ;
      RECT 12.735000  0.890000 13.360000 1.220000 ;
      RECT 13.020000  0.255000 13.360000 0.890000 ;
      RECT 13.020000  1.220000 13.360000 2.465000 ;
      RECT 13.530000  0.085000 13.765000 0.900000 ;
      RECT 13.530000  1.465000 13.765000 2.635000 ;
      RECT 14.435000  0.085000 14.695000 0.900000 ;
      RECT 14.435000  1.465000 14.695000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.615000  0.425000  4.785000 0.595000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.530000  0.425000  6.700000 0.595000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.100000  1.445000  7.270000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.510000  1.785000  7.680000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.100000  1.785000 10.270000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.520000  1.445000 10.690000 1.615000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.980000  1.785000 11.150000 1.955000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 12.650000  1.785000 12.820000 1.955000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.110000  0.765000 13.280000 0.935000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000 10.330000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000 10.750000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 13.340000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.555000 0.395000  6.760000 0.580000 ;
      RECT  4.555000 0.580000  4.845000 0.625000 ;
      RECT  6.470000 0.580000  6.760000 0.625000 ;
      RECT  7.040000 1.415000  7.330000 1.460000 ;
      RECT  7.040000 1.600000  7.330000 1.645000 ;
      RECT  7.450000 1.755000  7.740000 1.800000 ;
      RECT  7.450000 1.940000  7.740000 1.985000 ;
      RECT 10.040000 1.755000 10.330000 1.800000 ;
      RECT 10.040000 1.940000 10.330000 1.985000 ;
      RECT 10.460000 1.415000 10.750000 1.460000 ;
      RECT 10.460000 1.600000 10.750000 1.645000 ;
      RECT 10.920000 1.755000 11.210000 1.800000 ;
      RECT 10.920000 1.800000 12.880000 1.940000 ;
      RECT 10.920000 1.940000 11.210000 1.985000 ;
      RECT 12.590000 1.755000 12.880000 1.800000 ;
      RECT 12.590000 1.940000 12.880000 1.985000 ;
      RECT 13.050000 0.735000 13.340000 0.780000 ;
      RECT 13.050000 0.920000 13.340000 0.965000 ;
  END
END sky130_fd_sc_hd__sedfxbp_2
MACRO sky130_fd_sc_hd__sedfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.26000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.525000 0.255000 13.855000 2.420000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.700000 1.065000 12.145000 1.410000 ;
        RECT 11.700000 1.410000 12.030000 2.465000 ;
        RECT 11.815000 0.255000 12.145000 1.065000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 1.105000 6.215000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.105000 5.250000 1.615000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000  4.885000 1.435000 ;
        RECT -0.190000 1.435000 14.450000 2.910000 ;
        RECT  7.200000 1.305000 14.450000 1.435000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.595000  0.255000  4.795000 0.645000 ;
      RECT  4.595000  0.645000  4.855000 0.825000 ;
      RECT  4.635000  2.210000  4.965000 2.465000 ;
      RECT  4.685000  0.825000  4.855000 1.785000 ;
      RECT  4.685000  1.785000  4.965000 2.210000 ;
      RECT  4.965000  0.255000  5.590000 0.515000 ;
      RECT  5.155000  1.835000  6.585000 2.005000 ;
      RECT  5.155000  2.005000  5.495000 2.465000 ;
      RECT  5.260000  0.515000  5.590000 0.935000 ;
      RECT  5.420000  0.935000  5.590000 1.835000 ;
      RECT  5.665000  2.175000  6.010000 2.635000 ;
      RECT  5.760000  0.085000  6.010000 0.905000 ;
      RECT  6.385000  1.355000  6.585000 1.835000 ;
      RECT  6.515000  0.255000  7.135000 0.565000 ;
      RECT  6.515000  0.565000  6.925000 1.185000 ;
      RECT  6.675000  2.150000  7.005000 2.465000 ;
      RECT  6.755000  1.185000  6.925000 1.865000 ;
      RECT  6.755000  1.865000  7.005000 2.150000 ;
      RECT  7.095000  1.125000  7.280000 1.720000 ;
      RECT  7.115000  0.735000  7.620000 0.955000 ;
      RECT  7.215000  2.175000  8.255000 2.375000 ;
      RECT  7.305000  0.255000  7.980000 0.565000 ;
      RECT  7.450000  0.955000  7.620000 1.655000 ;
      RECT  7.450000  1.655000  7.915000 2.005000 ;
      RECT  7.810000  0.565000  7.980000 1.315000 ;
      RECT  7.810000  1.315000  8.660000 1.485000 ;
      RECT  8.085000  1.485000  8.660000 1.575000 ;
      RECT  8.085000  1.575000  8.255000 2.175000 ;
      RECT  8.170000  0.765000  9.235000 1.045000 ;
      RECT  8.170000  1.045000  9.745000 1.065000 ;
      RECT  8.170000  1.065000  8.370000 1.095000 ;
      RECT  8.245000  0.085000  8.640000 0.560000 ;
      RECT  8.425000  1.835000  8.660000 2.635000 ;
      RECT  8.490000  1.245000  8.660000 1.315000 ;
      RECT  8.830000  0.255000  9.235000 0.765000 ;
      RECT  8.830000  1.065000  9.745000 1.375000 ;
      RECT  8.830000  1.375000  9.160000 2.465000 ;
      RECT  9.370000  2.105000  9.660000 2.635000 ;
      RECT  9.465000  0.085000  9.740000 0.615000 ;
      RECT 10.090000  1.245000 10.280000 1.965000 ;
      RECT 10.225000  2.165000 11.190000 2.355000 ;
      RECT 10.305000  0.705000 10.770000 1.035000 ;
      RECT 10.325000  0.330000 11.190000 0.535000 ;
      RECT 10.450000  1.035000 10.770000 1.995000 ;
      RECT 10.940000  0.535000 11.190000 2.165000 ;
      RECT 11.360000  1.495000 11.530000 2.635000 ;
      RECT 11.395000  0.085000 11.645000 0.900000 ;
      RECT 12.200000  1.575000 12.430000 2.010000 ;
      RECT 12.315000  0.890000 12.940000 1.220000 ;
      RECT 12.600000  0.255000 12.940000 0.890000 ;
      RECT 12.600000  1.220000 12.940000 2.465000 ;
      RECT 13.110000  0.085000 13.355000 0.900000 ;
      RECT 13.110000  1.465000 13.355000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.615000  0.425000  4.785000 0.595000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.530000  0.425000  6.700000 0.595000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.100000  1.445000  7.270000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.510000  1.785000  7.680000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.100000  1.785000 10.270000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.520000  1.445000 10.690000 1.615000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 10.980000  1.785000 11.150000 1.955000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.230000  1.785000 12.400000 1.955000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 12.690000  0.765000 12.860000 0.935000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000 10.330000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000 10.750000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 12.920000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.555000 0.395000  6.760000 0.580000 ;
      RECT  4.555000 0.580000  4.845000 0.625000 ;
      RECT  6.470000 0.580000  6.760000 0.625000 ;
      RECT  7.040000 1.415000  7.330000 1.460000 ;
      RECT  7.040000 1.600000  7.330000 1.645000 ;
      RECT  7.450000 1.755000  7.740000 1.800000 ;
      RECT  7.450000 1.940000  7.740000 1.985000 ;
      RECT 10.040000 1.755000 10.330000 1.800000 ;
      RECT 10.040000 1.940000 10.330000 1.985000 ;
      RECT 10.460000 1.415000 10.750000 1.460000 ;
      RECT 10.460000 1.600000 10.750000 1.645000 ;
      RECT 10.920000 1.755000 11.210000 1.800000 ;
      RECT 10.920000 1.800000 12.460000 1.940000 ;
      RECT 10.920000 1.940000 11.210000 1.985000 ;
      RECT 12.170000 1.755000 12.460000 1.800000 ;
      RECT 12.170000 1.940000 12.460000 1.985000 ;
      RECT 12.630000 0.735000 12.920000 0.780000 ;
      RECT 12.630000 0.920000 12.920000 0.965000 ;
  END
END sky130_fd_sc_hd__sedfxbp_1
MACRO sky130_fd_sc_hd__nand4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.330000 1.615000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.010000 1.075000 3.100000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.360000 1.075000 4.450000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.620000 1.075000 5.430000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.635000 1.785000 0.825000 ;
        RECT 1.455000 1.445000 4.865000 1.665000 ;
        RECT 1.455000 1.665000 1.785000 2.465000 ;
        RECT 1.550000 0.825000 1.785000 1.445000 ;
        RECT 2.295000 1.665000 2.625000 2.465000 ;
        RECT 3.605000 1.665000 3.935000 2.465000 ;
        RECT 4.535000 1.665000 4.865000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.090000  0.255000 0.345000 0.635000 ;
      RECT 0.090000  0.635000 0.670000 0.805000 ;
      RECT 0.090000  1.915000 0.670000 2.085000 ;
      RECT 0.090000  2.085000 0.345000 2.465000 ;
      RECT 0.500000  0.805000 0.670000 1.075000 ;
      RECT 0.500000  1.075000 1.380000 1.245000 ;
      RECT 0.500000  1.245000 0.670000 1.915000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.255000 1.285000 2.635000 ;
      RECT 1.035000  0.255000 2.125000 0.465000 ;
      RECT 1.035000  0.465000 1.285000 0.905000 ;
      RECT 1.035000  1.445000 1.285000 2.255000 ;
      RECT 1.955000  0.465000 2.125000 0.635000 ;
      RECT 1.955000  0.635000 3.045000 0.905000 ;
      RECT 1.955000  1.835000 2.125000 2.635000 ;
      RECT 2.295000  0.255000 3.985000 0.465000 ;
      RECT 2.795000  1.835000 3.435000 2.635000 ;
      RECT 3.235000  0.635000 4.455000 0.715000 ;
      RECT 3.235000  0.715000 5.340000 0.905000 ;
      RECT 4.105000  1.835000 4.365000 2.635000 ;
      RECT 4.155000  0.255000 4.415000 0.615000 ;
      RECT 4.155000  0.615000 4.455000 0.635000 ;
      RECT 4.665000  0.085000 4.835000 0.545000 ;
      RECT 5.005000  0.255000 5.340000 0.715000 ;
      RECT 5.035000  1.495000 5.430000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4b_2
MACRO sky130_fd_sc_hd__nand4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.930000 1.075000 4.590000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.790000 1.075000 6.510000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.015000 1.075000 8.655000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.635000 2.640000 0.905000 ;
        RECT 1.455000 1.445000 8.185000 1.665000 ;
        RECT 1.455000 1.665000 1.785000 2.465000 ;
        RECT 2.295000 1.665000 2.625000 2.465000 ;
        RECT 2.375000 0.905000 2.640000 1.445000 ;
        RECT 3.135000 1.665000 3.465000 2.465000 ;
        RECT 3.975000 1.665000 4.305000 2.465000 ;
        RECT 5.335000 1.665000 5.665000 2.465000 ;
        RECT 6.175000 1.665000 6.505000 2.465000 ;
        RECT 7.015000 1.665000 7.345000 2.465000 ;
        RECT 7.855000 1.665000 8.185000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 0.805000 0.905000 ;
      RECT 0.090000  1.495000 0.805000 1.665000 ;
      RECT 0.090000  1.665000 0.425000 2.465000 ;
      RECT 0.595000  0.085000 0.845000 0.545000 ;
      RECT 0.595000  1.835000 1.285000 2.635000 ;
      RECT 0.610000  0.905000 0.805000 1.075000 ;
      RECT 0.610000  1.075000 2.205000 1.275000 ;
      RECT 0.610000  1.275000 0.805000 1.495000 ;
      RECT 0.995000  1.495000 1.285000 1.835000 ;
      RECT 1.035000  0.255000 4.725000 0.465000 ;
      RECT 1.035000  0.465000 1.285000 0.905000 ;
      RECT 1.955000  1.835000 2.125000 2.635000 ;
      RECT 2.795000  1.835000 2.965000 2.635000 ;
      RECT 3.135000  0.635000 6.505000 0.905000 ;
      RECT 3.635000  1.835000 3.805000 2.635000 ;
      RECT 4.475000  1.835000 5.165000 2.635000 ;
      RECT 4.915000  0.255000 6.925000 0.465000 ;
      RECT 5.835000  1.835000 6.005000 2.635000 ;
      RECT 6.675000  0.465000 6.925000 0.735000 ;
      RECT 6.675000  0.735000 8.610000 0.905000 ;
      RECT 6.675000  1.835000 6.845000 2.635000 ;
      RECT 7.095000  0.085000 7.265000 0.545000 ;
      RECT 7.435000  0.255000 7.765000 0.735000 ;
      RECT 7.515000  1.835000 7.685000 2.635000 ;
      RECT 7.935000  0.085000 8.105000 0.545000 ;
      RECT 8.275000  0.255000 8.610000 0.735000 ;
      RECT 8.355000  1.445000 8.610000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4b_4
MACRO sky130_fd_sc_hd__nand4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 0.765000 2.185000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 0.765000 1.755000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 0.995000 1.235000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.887500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.130000 1.495000 3.135000 1.665000 ;
        RECT 1.130000 1.665000 1.460000 2.465000 ;
        RECT 2.085000 1.665000 2.415000 2.465000 ;
        RECT 2.695000 0.255000 3.135000 0.825000 ;
        RECT 2.925000 0.825000 3.135000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.445000 0.475000 0.655000 ;
      RECT 0.085000  0.655000 1.335000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.595000 ;
      RECT 0.085000  1.595000 0.510000 1.925000 ;
      RECT 0.655000  0.085000 0.985000 0.485000 ;
      RECT 0.710000  1.495000 0.960000 2.635000 ;
      RECT 1.155000  0.425000 2.525000 0.595000 ;
      RECT 1.155000  0.595000 1.335000 0.655000 ;
      RECT 1.630000  1.835000 1.915000 2.635000 ;
      RECT 2.355000  0.595000 2.525000 0.995000 ;
      RECT 2.355000  0.995000 2.755000 1.325000 ;
      RECT 2.705000  1.835000 2.920000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4b_1
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.545000 1.755000 2.465000 ;
        RECT 1.005000 1.025000 1.755000 1.545000 ;
      LAYER mcon ;
        RECT 0.145000 2.125000 0.315000 2.295000 ;
        RECT 0.605000 2.125000 0.775000 2.295000 ;
        RECT 1.065000 2.125000 1.235000 2.295000 ;
        RECT 1.525000 2.125000 1.695000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 1.770000 2.340000 ;
        RECT 0.085000 2.080000 1.755000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.085000 1.755000 0.855000 ;
      RECT 0.085000  0.855000 0.835000 1.375000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_4
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_3
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_3 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.545000 1.295000 2.465000 ;
        RECT 0.775000 1.005000 1.295000 1.545000 ;
      LAYER mcon ;
        RECT 0.145000 2.125000 0.315000 2.295000 ;
        RECT 0.605000 2.125000 0.775000 2.295000 ;
        RECT 1.065000 2.125000 1.235000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 1.310000 2.340000 ;
        RECT 0.085000 2.080000 1.295000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.085000  0.085000 1.295000 0.835000 ;
      RECT 0.085000  0.835000 0.605000 1.375000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_3
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.545000 3.595000 2.465000 ;
        RECT 1.905000 1.025000 3.595000 1.545000 ;
      LAYER mcon ;
        RECT 0.145000 2.125000 0.315000 2.295000 ;
        RECT 0.605000 2.125000 0.775000 2.295000 ;
        RECT 1.065000 2.125000 1.235000 2.295000 ;
        RECT 1.525000 2.125000 1.695000 2.295000 ;
        RECT 1.985000 2.125000 2.155000 2.295000 ;
        RECT 2.445000 2.125000 2.615000 2.295000 ;
        RECT 2.905000 2.125000 3.075000 2.295000 ;
        RECT 3.365000 2.125000 3.535000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 3.610000 2.340000 ;
        RECT 0.085000 2.080000 3.595000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 3.595000 0.855000 ;
      RECT 0.085000  0.855000 1.735000 1.375000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_8
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.545000 5.430000 2.465000 ;
        RECT 2.835000 1.025000 5.430000 1.545000 ;
      LAYER mcon ;
        RECT 0.145000 2.125000 0.315000 2.295000 ;
        RECT 0.605000 2.125000 0.775000 2.295000 ;
        RECT 1.065000 2.125000 1.235000 2.295000 ;
        RECT 1.525000 2.125000 1.695000 2.295000 ;
        RECT 1.985000 2.125000 2.155000 2.295000 ;
        RECT 2.445000 2.125000 2.615000 2.295000 ;
        RECT 2.905000 2.125000 3.075000 2.295000 ;
        RECT 3.365000 2.125000 3.535000 2.295000 ;
        RECT 3.825000 2.125000 3.995000 2.295000 ;
        RECT 4.285000 2.125000 4.455000 2.295000 ;
        RECT 4.745000 2.125000 4.915000 2.295000 ;
        RECT 5.205000 2.125000 5.375000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 5.450000 2.340000 ;
        RECT 0.085000 2.080000 5.435000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.085000 5.430000 0.855000 ;
      RECT 0.085000  0.855000 2.665000 1.375000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_12
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.545000 2.675000 2.465000 ;
        RECT 1.465000 1.025000 2.675000 1.545000 ;
      LAYER mcon ;
        RECT 0.145000 2.125000 0.315000 2.295000 ;
        RECT 0.605000 2.125000 0.775000 2.295000 ;
        RECT 1.065000 2.125000 1.235000 2.295000 ;
        RECT 1.525000 2.125000 1.695000 2.295000 ;
        RECT 1.985000 2.125000 2.155000 2.295000 ;
        RECT 2.445000 2.125000 2.615000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 2.690000 2.340000 ;
        RECT 0.085000 2.080000 2.675000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.085000 2.675000 0.855000 ;
      RECT 0.085000  0.855000 1.295000 1.375000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_6
MACRO sky130_fd_sc_hd__mux2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 0.255000 2.265000 1.415000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.615000 0.815000 1.785000 1.615000 ;
        RECT 1.615000 1.615000 2.625000 1.785000 ;
        RECT 2.435000 0.255000 2.625000 1.615000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 0.995000 1.105000 1.325000 ;
        RECT 0.935000 1.325000 1.105000 2.295000 ;
        RECT 0.935000 2.295000 2.965000 2.465000 ;
        RECT 2.795000 1.440000 3.545000 1.630000 ;
        RECT 2.795000 1.630000 2.965000 2.295000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.255000 0.345000 0.825000 ;
        RECT 0.090000 0.825000 0.260000 1.495000 ;
        RECT 0.090000 1.495000 0.425000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.420000 -0.085000 0.590000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.430000  0.995000 0.685000 1.325000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  0.655000 1.445000 0.825000 ;
      RECT 0.515000  0.825000 0.685000 0.995000 ;
      RECT 0.595000  1.495000 0.765000 2.635000 ;
      RECT 1.270000  0.255000 1.800000 0.620000 ;
      RECT 1.270000  0.620000 1.445000 0.655000 ;
      RECT 1.275000  0.825000 1.445000 1.955000 ;
      RECT 1.275000  1.955000 2.400000 2.125000 ;
      RECT 2.805000  0.085000 3.315000 0.620000 ;
      RECT 2.825000  0.895000 4.055000 1.065000 ;
      RECT 3.135000  1.875000 3.305000 2.635000 ;
      RECT 3.535000  0.290000 3.780000 0.895000 ;
      RECT 3.540000  1.875000 4.055000 2.285000 ;
      RECT 3.715000  1.065000 4.055000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__mux2_1
MACRO sky130_fd_sc_hd__mux2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 0.995000 1.750000 1.615000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 0.995000 2.435000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.740000 1.325000 ;
        RECT 0.570000 0.635000 2.850000 0.805000 ;
        RECT 0.570000 0.805000 0.740000 0.995000 ;
        RECT 2.680000 0.805000 2.850000 0.995000 ;
        RECT 2.680000 0.995000 3.395000 1.325000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.915000 0.255000 4.085000 0.635000 ;
        RECT 3.915000 0.635000 5.430000 0.805000 ;
        RECT 3.915000 1.575000 5.430000 1.745000 ;
        RECT 3.915000 1.745000 4.085000 2.465000 ;
        RECT 4.755000 0.255000 4.925000 0.635000 ;
        RECT 4.755000 1.745000 4.925000 2.465000 ;
        RECT 5.200000 0.805000 5.430000 1.575000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.090000  0.295000 0.345000 0.625000 ;
      RECT 0.090000  0.625000 0.260000 1.495000 ;
      RECT 0.090000  1.495000 1.080000 1.665000 ;
      RECT 0.090000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  1.835000 0.820000 2.635000 ;
      RECT 0.910000  0.995000 1.080000 1.495000 ;
      RECT 0.990000  1.935000 1.340000 2.275000 ;
      RECT 0.990000  2.275000 2.770000 2.445000 ;
      RECT 1.530000  1.935000 3.245000 2.105000 ;
      RECT 1.975000  0.295000 3.230000 0.465000 ;
      RECT 1.980000  1.595000 3.735000 1.765000 ;
      RECT 3.060000  0.465000 3.230000 0.655000 ;
      RECT 3.060000  0.655000 3.735000 0.825000 ;
      RECT 3.075000  2.105000 3.245000 2.465000 ;
      RECT 3.415000  0.085000 3.745000 0.465000 ;
      RECT 3.415000  2.255000 3.745000 2.635000 ;
      RECT 3.565000  0.825000 3.735000 1.075000 ;
      RECT 3.565000  1.075000 5.030000 1.245000 ;
      RECT 3.565000  1.245000 3.735000 1.595000 ;
      RECT 3.565000  1.765000 3.735000 1.785000 ;
      RECT 4.255000  0.085000 4.585000 0.465000 ;
      RECT 4.255000  1.915000 4.585000 2.635000 ;
      RECT 5.095000  0.085000 5.425000 0.465000 ;
      RECT 5.095000  1.915000 5.425000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__mux2_4
MACRO sky130_fd_sc_hd__mux2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.815000 0.765000 2.445000 1.280000 ;
        RECT 2.275000 1.280000 2.445000 1.315000 ;
        RECT 2.275000 1.315000 3.090000 1.625000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.625000 0.735000 3.090000 1.025000 ;
        RECT 2.900000 0.420000 3.090000 0.735000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.360000 0.755000 3.550000 1.625000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.765000 0.750000 ;
        RECT 0.515000 0.750000 0.685000 1.595000 ;
        RECT 0.515000 1.595000 0.825000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.885000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.855000  0.995000 1.165000 1.325000 ;
      RECT 0.935000  0.085000 1.265000 0.465000 ;
      RECT 0.995000  0.635000 1.605000 0.805000 ;
      RECT 0.995000  0.805000 1.165000 0.995000 ;
      RECT 0.995000  1.325000 1.165000 1.835000 ;
      RECT 0.995000  1.835000 1.655000 2.005000 ;
      RECT 1.025000  2.175000 1.315000 2.635000 ;
      RECT 1.335000  0.995000 1.505000 1.495000 ;
      RECT 1.335000  1.495000 1.995000 1.665000 ;
      RECT 1.435000  0.295000 2.730000 0.465000 ;
      RECT 1.435000  0.465000 1.605000 0.635000 ;
      RECT 1.485000  2.005000 1.655000 2.255000 ;
      RECT 1.485000  2.255000 2.795000 2.425000 ;
      RECT 1.825000  1.665000 1.995000 1.835000 ;
      RECT 1.825000  1.835000 4.050000 2.005000 ;
      RECT 3.325000  2.175000 3.545000 2.635000 ;
      RECT 3.350000  0.085000 3.550000 0.585000 ;
      RECT 3.715000  2.005000 4.050000 2.465000 ;
      RECT 3.720000  0.255000 4.050000 1.835000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__mux2_2
MACRO sky130_fd_sc_hd__mux2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.180000 0.645000 6.895000 0.815000 ;
        RECT 5.180000 0.815000 5.350000 1.325000 ;
        RECT 5.305000 0.425000 5.890000 0.645000 ;
        RECT 6.725000 0.815000 6.895000 0.995000 ;
        RECT 6.725000 0.995000 7.195000 1.165000 ;
        RECT 7.025000 1.165000 7.195000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.290000 1.105000 4.475000 1.275000 ;
        RECT 4.305000 0.995000 4.475000 1.105000 ;
        RECT 4.305000 1.275000 4.475000 1.325000 ;
      LAYER mcon ;
        RECT 4.290000 1.105000 4.460000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.960000 0.995000 8.245000 1.325000 ;
      LAYER mcon ;
        RECT 7.960000 1.105000 8.130000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.230000 1.075000 4.520000 1.120000 ;
        RECT 4.230000 1.120000 8.190000 1.260000 ;
        RECT 4.230000 1.260000 4.520000 1.305000 ;
        RECT 7.900000 1.075000 8.190000 1.120000 ;
        RECT 7.900000 1.260000 8.190000 1.305000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.739500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.795000 0.995000 3.965000 1.495000 ;
        RECT 3.795000 1.495000 6.035000 1.665000 ;
        RECT 5.670000 0.995000 6.035000 1.495000 ;
      LAYER mcon ;
        RECT 5.670000 1.445000 5.840000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.215000 0.995000 9.510000 1.615000 ;
      LAYER mcon ;
        RECT 9.340000 1.445000 9.510000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.610000 1.415000 5.900000 1.460000 ;
        RECT 5.610000 1.460000 9.570000 1.600000 ;
        RECT 5.610000 1.600000 5.900000 1.645000 ;
        RECT 9.280000 1.415000 9.570000 1.460000 ;
        RECT 9.280000 1.600000 9.570000 1.645000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.255000 0.765000 0.635000 ;
        RECT 0.595000 0.635000 3.285000 0.805000 ;
        RECT 0.595000 0.805000 0.815000 1.575000 ;
        RECT 0.595000 1.575000 3.285000 1.745000 ;
        RECT 0.595000 1.745000 0.765000 2.465000 ;
        RECT 1.435000 0.295000 1.605000 0.635000 ;
        RECT 1.435000 1.745000 1.605000 2.465000 ;
        RECT 2.275000 0.255000 2.445000 0.635000 ;
        RECT 2.275000 1.745000 2.445000 2.465000 ;
        RECT 3.115000 0.295000 3.285000 0.635000 ;
        RECT 3.115000 1.745000 3.285000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.465000 ;
      RECT 0.090000  1.915000 0.425000 2.635000 ;
      RECT 0.935000  0.085000 1.265000 0.465000 ;
      RECT 0.935000  1.915000 1.265000 2.635000 ;
      RECT 0.985000  1.075000 3.625000 1.245000 ;
      RECT 1.775000  0.085000 2.105000 0.465000 ;
      RECT 1.775000  1.915000 2.105000 2.635000 ;
      RECT 2.615000  0.085000 2.945000 0.465000 ;
      RECT 2.615000  1.915000 2.945000 2.635000 ;
      RECT 3.455000  0.085000 3.785000 0.465000 ;
      RECT 3.455000  0.635000 4.920000 0.805000 ;
      RECT 3.455000  0.805000 3.625000 1.075000 ;
      RECT 3.455000  1.245000 3.625000 1.835000 ;
      RECT 3.455000  1.835000 8.225000 2.005000 ;
      RECT 3.455000  2.255000 3.785000 2.635000 ;
      RECT 3.955000  0.295000 5.125000 0.465000 ;
      RECT 3.955000  2.255000 5.905000 2.425000 ;
      RECT 4.750000  0.805000 4.920000 0.935000 ;
      RECT 6.060000  0.085000 6.390000 0.465000 ;
      RECT 6.075000  2.175000 6.245000 2.635000 ;
      RECT 6.345000  0.995000 6.515000 1.495000 ;
      RECT 6.345000  1.495000 8.855000 1.665000 ;
      RECT 6.480000  2.255000 8.645000 2.425000 ;
      RECT 6.575000  0.295000 7.865000 0.465000 ;
      RECT 7.115000  0.635000 7.670000 0.805000 ;
      RECT 7.500000  0.805000 7.670000 0.935000 ;
      RECT 8.685000  0.645000 9.485000 0.815000 ;
      RECT 8.685000  0.815000 8.855000 1.495000 ;
      RECT 8.685000  1.665000 8.855000 1.915000 ;
      RECT 8.685000  1.915000 9.485000 2.085000 ;
      RECT 8.815000  0.085000 9.145000 0.465000 ;
      RECT 8.815000  2.255000 9.145000 2.635000 ;
      RECT 9.315000  0.295000 9.485000 0.645000 ;
      RECT 9.315000  1.795000 9.485000 1.915000 ;
      RECT 9.315000  2.085000 9.485000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 4.750000  0.765000 4.920000 0.935000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.500000  0.765000 7.670000 0.935000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 4.690000 0.735000 4.980000 0.780000 ;
      RECT 4.690000 0.780000 7.730000 0.920000 ;
      RECT 4.690000 0.920000 4.980000 0.965000 ;
      RECT 7.440000 0.735000 7.730000 0.780000 ;
      RECT 7.440000 0.920000 7.730000 0.965000 ;
  END
END sky130_fd_sc_hd__mux2_8
MACRO sky130_fd_sc_hd__a311oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.000000 0.995000 3.115000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 0.995000 1.805000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.995000 0.800000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 0.995000 4.055000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.730000 1.075000 5.410000 1.295000 ;
        RECT 5.175000 1.295000 5.410000 1.625000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.141000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 0.655000 5.345000 0.825000 ;
        RECT 3.235000 0.255000 3.405000 0.655000 ;
        RECT 4.085000 0.255000 4.255000 0.655000 ;
        RECT 4.260000 0.825000 4.475000 1.510000 ;
        RECT 4.260000 1.510000 4.990000 1.575000 ;
        RECT 4.260000 1.575000 5.005000 1.680000 ;
        RECT 4.660000 1.680000 5.005000 1.745000 ;
        RECT 4.660000 1.745000 4.990000 1.915000 ;
        RECT 4.660000 1.915000 5.005000 2.085000 ;
        RECT 5.175000 0.255000 5.345000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.095000  1.495000 0.345000 2.635000 ;
      RECT 0.175000  0.255000 0.345000 0.655000 ;
      RECT 0.175000  0.655000 2.105000 0.825000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.595000  1.575000 3.915000 1.745000 ;
      RECT 0.595000  1.745000 0.765000 2.465000 ;
      RECT 0.935000  1.915000 1.265000 2.635000 ;
      RECT 1.015000  0.255000 1.185000 0.655000 ;
      RECT 1.355000  0.305000 3.045000 0.475000 ;
      RECT 1.435000  1.745000 1.605000 2.465000 ;
      RECT 1.785000  1.915000 2.135000 2.635000 ;
      RECT 2.305000  1.745000 2.475000 2.465000 ;
      RECT 2.645000  1.915000 2.975000 2.635000 ;
      RECT 3.145000  2.255000 5.345000 2.425000 ;
      RECT 3.585000  0.085000 3.915000 0.465000 ;
      RECT 3.585000  1.745000 3.915000 2.085000 ;
      RECT 4.110000  1.915000 4.440000 2.255000 ;
      RECT 4.110000  2.425000 4.440000 2.465000 ;
      RECT 4.675000  0.085000 5.005000 0.465000 ;
      RECT 5.175000  1.795000 5.345000 2.255000 ;
      RECT 5.175000  2.425000 5.345000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__a311oi_2
MACRO sky130_fd_sc_hd__a311oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.995000 5.420000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.995000 3.550000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.995000 1.735000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.670000 0.995000 6.855000 1.630000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.935000 0.995000 9.530000 1.325000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.898500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.975000 0.635000 9.485000 0.805000 ;
        RECT 6.575000 0.255000 6.745000 0.635000 ;
        RECT 7.415000 0.255000 7.585000 0.635000 ;
        RECT 7.415000 0.805000 7.735000 1.545000 ;
        RECT 7.415000 1.545000 9.145000 1.715000 ;
        RECT 7.415000 1.715000 7.735000 1.975000 ;
        RECT 7.975000 1.530000 8.305000 1.545000 ;
        RECT 7.975000 1.715000 8.305000 2.085000 ;
        RECT 8.475000 0.255000 8.645000 0.635000 ;
        RECT 8.815000 1.715000 9.145000 2.085000 ;
        RECT 9.315000 0.255000 9.485000 0.635000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.095000  1.575000 0.425000 2.635000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 3.785000 0.805000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.595000  1.495000 4.965000 1.665000 ;
      RECT 0.595000  1.665000 0.765000 2.465000 ;
      RECT 0.935000  1.915000 1.265000 2.635000 ;
      RECT 1.015000  0.255000 1.185000 0.635000 ;
      RECT 1.355000  0.085000 1.685000 0.465000 ;
      RECT 1.435000  1.665000 1.605000 2.465000 ;
      RECT 1.775000  1.915000 2.105000 2.635000 ;
      RECT 1.855000  0.255000 2.025000 0.635000 ;
      RECT 2.195000  0.295000 5.565000 0.465000 ;
      RECT 2.275000  1.665000 2.445000 2.465000 ;
      RECT 2.615000  1.915000 2.945000 2.635000 ;
      RECT 3.115000  1.665000 3.285000 2.465000 ;
      RECT 3.455000  1.915000 3.785000 2.635000 ;
      RECT 3.955000  1.665000 4.125000 2.465000 ;
      RECT 4.295000  1.915000 4.625000 2.635000 ;
      RECT 4.795000  1.665000 4.965000 1.915000 ;
      RECT 4.795000  1.915000 7.245000 2.085000 ;
      RECT 4.795000  2.085000 4.965000 2.465000 ;
      RECT 5.135000  2.255000 5.465000 2.635000 ;
      RECT 5.655000  2.255000 9.565000 2.425000 ;
      RECT 6.075000  0.085000 6.405000 0.465000 ;
      RECT 6.915000  0.085000 7.245000 0.465000 ;
      RECT 7.975000  0.085000 8.305000 0.465000 ;
      RECT 8.815000  0.085000 9.145000 0.465000 ;
      RECT 9.315000  1.835000 9.565000 2.255000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__a311oi_4
MACRO sky130_fd_sc_hd__a311oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 0.265000 1.365000 0.660000 ;
        RECT 1.195000 0.660000 1.365000 0.995000 ;
        RECT 1.195000 0.995000 1.455000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.600000 0.265000 0.795000 0.995000 ;
        RECT 0.600000 0.995000 1.025000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.420000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.710000 0.995000 1.935000 1.835000 ;
        RECT 1.710000 1.835000 2.230000 2.005000 ;
        RECT 1.950000 2.005000 2.230000 2.355000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.995000 2.685000 1.325000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.659750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 0.255000 1.705000 0.655000 ;
        RECT 1.535000 0.655000 2.650000 0.825000 ;
        RECT 2.105000 0.825000 2.275000 1.495000 ;
        RECT 2.105000 1.495000 2.650000 1.665000 ;
        RECT 2.405000 0.295000 2.650000 0.655000 ;
        RECT 2.410000 1.665000 2.650000 2.335000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.805000 ;
      RECT 0.095000  1.495000 0.425000 2.635000 ;
      RECT 0.600000  1.575000 1.540000 1.745000 ;
      RECT 0.600000  1.745000 0.770000 2.305000 ;
      RECT 0.940000  1.915000 1.200000 2.635000 ;
      RECT 1.370000  1.745000 1.540000 2.175000 ;
      RECT 1.370000  2.175000 1.700000 2.345000 ;
      RECT 1.905000  0.085000 2.235000 0.485000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a311oi_1
MACRO sky130_fd_sc_hd__probe_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__probe_p_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.240000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1.250000 0.560000 4.270000 2.160000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.095000  1.445000 1.595000 1.615000 ;
      RECT 0.095000  1.615000 0.425000 2.465000 ;
      RECT 0.175000  0.255000 0.345000 0.735000 ;
      RECT 0.175000  0.735000 1.595000 0.905000 ;
      RECT 0.515000  0.085000 0.845000 0.565000 ;
      RECT 0.595000  1.835000 0.765000 2.635000 ;
      RECT 0.935000  1.615000 1.265000 2.465000 ;
      RECT 1.015000  0.260000 1.185000 0.735000 ;
      RECT 1.355000  0.085000 1.685000 0.565000 ;
      RECT 1.420000  0.905000 1.595000 1.075000 ;
      RECT 1.420000  1.075000 4.045000 1.245000 ;
      RECT 1.420000  1.245000 1.595000 1.445000 ;
      RECT 1.435000  1.835000 1.605000 2.635000 ;
      RECT 1.855000  0.255000 2.025000 0.735000 ;
      RECT 1.855000  0.735000 4.545000 0.905000 ;
      RECT 1.855000  1.445000 4.545000 1.615000 ;
      RECT 1.855000  1.615000 2.025000 2.465000 ;
      RECT 2.195000  0.085000 2.525000 0.565000 ;
      RECT 2.195000  1.835000 2.525000 2.635000 ;
      RECT 2.695000  0.255000 2.865000 0.735000 ;
      RECT 2.695000  1.615000 2.865000 2.465000 ;
      RECT 3.035000  0.085000 3.365000 0.565000 ;
      RECT 3.035000  1.835000 3.365000 2.635000 ;
      RECT 3.535000  0.255000 3.705000 0.735000 ;
      RECT 3.535000  1.615000 3.705000 2.465000 ;
      RECT 3.875000  0.085000 4.205000 0.565000 ;
      RECT 3.875000  1.835000 4.205000 2.635000 ;
      RECT 4.290000  0.905000 4.545000 1.055000 ;
      RECT 4.290000  1.055000 4.885000 1.315000 ;
      RECT 4.290000  1.315000 4.545000 1.445000 ;
      RECT 4.375000  0.255000 4.545000 0.735000 ;
      RECT 4.375000  1.615000 4.545000 2.465000 ;
      RECT 4.715000  0.085000 5.045000 0.885000 ;
      RECT 4.715000  1.485000 5.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.320000  1.105000 4.490000 1.275000 ;
      RECT 4.680000  1.105000 4.850000 1.275000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
    LAYER met1 ;
      RECT 3.465000 1.060000 4.105000 1.075000 ;
      RECT 3.465000 1.075000 4.910000 1.305000 ;
      RECT 3.465000 1.305000 4.105000 1.320000 ;
    LAYER met2 ;
      RECT 3.445000 1.005000 4.125000 1.375000 ;
    LAYER met3 ;
      RECT 3.395000 1.025000 4.175000 1.355000 ;
    LAYER met4 ;
      RECT 1.370000 0.680000 4.150000 1.860000 ;
    LAYER via ;
      RECT 3.495000 1.060000 3.755000 1.320000 ;
      RECT 3.815000 1.060000 4.075000 1.320000 ;
    LAYER via2 ;
      RECT 3.445000 1.050000 3.725000 1.330000 ;
      RECT 3.845000 1.050000 4.125000 1.330000 ;
    LAYER via3 ;
      RECT 3.425000 1.030000 3.745000 1.350000 ;
      RECT 3.825000 1.030000 4.145000 1.350000 ;
    LAYER via4 ;
      RECT 2.970000 0.680000 4.150000 1.860000 ;
  END
END sky130_fd_sc_hd__probe_p_8
MACRO sky130_fd_sc_hd__xor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.075000 0.875000 1.275000 ;
        RECT 0.705000 1.275000 0.875000 1.445000 ;
        RECT 0.705000 1.445000 1.880000 1.615000 ;
        RECT 1.710000 1.075000 3.230000 1.275000 ;
        RECT 1.710000 1.275000 1.880000 1.445000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.075000 1.540000 1.275000 ;
      LAYER mcon ;
        RECT 1.065000 1.105000 1.235000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.420000 1.075000 4.090000 1.275000 ;
      LAYER mcon ;
        RECT 3.825000 1.105000 3.995000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.005000 1.075000 1.295000 1.120000 ;
        RECT 1.005000 1.120000 4.055000 1.260000 ;
        RECT 1.005000 1.260000 1.295000 1.305000 ;
        RECT 3.765000 1.075000 4.055000 1.120000 ;
        RECT 3.765000 1.260000 4.055000 1.305000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.656750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.625000 0.645000 3.955000 0.725000 ;
        RECT 3.625000 0.725000 5.895000 0.905000 ;
        RECT 4.985000 0.645000 5.315000 0.725000 ;
        RECT 5.025000 1.415000 5.895000 1.625000 ;
        RECT 5.025000 1.625000 5.275000 2.125000 ;
        RECT 5.485000 0.905000 5.895000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.120000  0.725000 1.700000 0.905000 ;
      RECT 0.120000  0.905000 0.290000 1.785000 ;
      RECT 0.120000  1.785000 2.220000 1.955000 ;
      RECT 0.120000  2.135000 0.400000 2.465000 ;
      RECT 0.145000  2.125000 0.315000 2.135000 ;
      RECT 0.190000  0.085000 0.360000 0.555000 ;
      RECT 0.530000  0.255000 0.860000 0.725000 ;
      RECT 0.570000  2.135000 0.820000 2.635000 ;
      RECT 0.990000  2.135000 1.240000 2.295000 ;
      RECT 0.990000  2.295000 2.080000 2.465000 ;
      RECT 1.030000  0.085000 1.200000 0.555000 ;
      RECT 1.065000  2.125000 1.235000 2.135000 ;
      RECT 1.370000  0.255000 1.700000 0.725000 ;
      RECT 1.410000  1.955000 1.660000 2.125000 ;
      RECT 1.830000  2.135000 2.080000 2.295000 ;
      RECT 1.870000  0.085000 2.040000 0.555000 ;
      RECT 2.050000  1.445000 4.785000 1.615000 ;
      RECT 2.050000  1.615000 2.220000 1.785000 ;
      RECT 2.285000  2.125000 2.600000 2.465000 ;
      RECT 2.310000  0.255000 2.640000 0.725000 ;
      RECT 2.310000  0.725000 3.400000 0.905000 ;
      RECT 2.390000  1.785000 4.855000 1.955000 ;
      RECT 2.390000  1.955000 2.600000 2.125000 ;
      RECT 2.770000  2.135000 3.020000 2.635000 ;
      RECT 2.810000  0.085000 2.980000 0.555000 ;
      RECT 3.150000  0.255000 4.380000 0.475000 ;
      RECT 3.150000  0.475000 3.400000 0.725000 ;
      RECT 3.190000  1.955000 3.440000 2.465000 ;
      RECT 3.610000  2.135000 3.915000 2.635000 ;
      RECT 4.085000  1.955000 4.855000 2.295000 ;
      RECT 4.085000  2.295000 5.695000 2.465000 ;
      RECT 4.615000  1.075000 5.275000 1.245000 ;
      RECT 4.615000  1.245000 4.785000 1.445000 ;
      RECT 4.645000  0.085000 4.815000 0.555000 ;
      RECT 5.445000  1.795000 5.695000 2.295000 ;
      RECT 5.485000  0.085000 5.655000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 0.085000 2.095000 0.375000 2.140000 ;
      RECT 0.085000 2.140000 1.295000 2.280000 ;
      RECT 0.085000 2.280000 0.375000 2.325000 ;
      RECT 1.005000 2.095000 1.295000 2.140000 ;
      RECT 1.005000 2.280000 1.295000 2.325000 ;
  END
END sky130_fd_sc_hd__xor2_2
MACRO sky130_fd_sc_hd__xor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.840000 1.075000 1.390000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.670000 1.445000 ;
        RECT 0.425000 1.445000 1.730000 1.615000 ;
        RECT 1.560000 1.075000 1.935000 1.245000 ;
        RECT 1.560000 1.245000 1.730000 1.445000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.800500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.720000 0.315000 2.675000 0.485000 ;
        RECT 2.505000 0.485000 2.675000 1.365000 ;
        RECT 2.505000 1.365000 3.135000 1.535000 ;
        RECT 2.815000 1.535000 3.135000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.655000 2.335000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.785000 ;
      RECT 0.085000  1.785000 0.465000 2.465000 ;
      RECT 0.135000  0.085000 0.465000 0.475000 ;
      RECT 0.635000  0.335000 0.805000 0.655000 ;
      RECT 0.975000  0.085000 1.305000 0.475000 ;
      RECT 1.055000  1.785000 1.225000 2.635000 ;
      RECT 1.395000  1.785000 2.635000 1.955000 ;
      RECT 1.395000  1.955000 1.725000 2.465000 ;
      RECT 1.895000  2.125000 2.065000 2.635000 ;
      RECT 2.105000  0.825000 2.335000 1.325000 ;
      RECT 2.235000  1.955000 2.635000 2.465000 ;
      RECT 2.845000  0.085000 3.135000 0.920000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__xor2_1
MACRO sky130_fd_sc_hd__xor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 2.800000 1.275000 ;
        RECT 2.630000 1.275000 2.800000 1.445000 ;
        RECT 2.630000 1.445000 6.165000 1.615000 ;
        RECT 5.995000 1.075000 7.370000 1.275000 ;
        RECT 5.995000 1.275000 6.165000 1.445000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.075000 5.000000 1.105000 ;
        RECT 2.970000 1.105000 5.740000 1.275000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.524450 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 0.645000 5.580000 0.905000 ;
        RECT 5.150000 0.905000 5.580000 0.935000 ;
      LAYER mcon ;
        RECT 5.205000 0.765000 5.375000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.850000 0.725000  8.630000 0.735000 ;
        RECT 7.850000 0.735000 10.035000 0.905000 ;
        RECT 7.850000 0.905000  8.305000 0.935000 ;
        RECT 7.880000 1.445000 10.035000 1.625000 ;
        RECT 7.880000 1.625000  9.010000 1.665000 ;
        RECT 7.880000 1.665000  8.170000 2.125000 ;
        RECT 8.300000 0.255000  8.630000 0.725000 ;
        RECT 8.760000 1.665000  9.010000 2.125000 ;
        RECT 9.140000 0.255000  9.470000 0.735000 ;
        RECT 9.600000 1.625000 10.035000 2.465000 ;
        RECT 9.735000 0.905000 10.035000 1.445000 ;
      LAYER mcon ;
        RECT 7.965000 0.765000 8.135000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.145000 0.735000 5.435000 0.780000 ;
        RECT 5.145000 0.780000 8.195000 0.920000 ;
        RECT 5.145000 0.920000 5.435000 0.965000 ;
        RECT 7.905000 0.735000 8.195000 0.780000 ;
        RECT 7.905000 0.920000 8.195000 0.965000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.085000  0.360000 0.565000 ;
      RECT 0.085000  0.735000  3.380000 0.905000 ;
      RECT 0.085000  0.905000  0.255000 1.445000 ;
      RECT 0.085000  1.445000  2.420000 1.615000 ;
      RECT 0.085000  1.785000  2.080000 2.005000 ;
      RECT 0.085000  2.005000  0.400000 2.465000 ;
      RECT 0.530000  0.255000  0.860000 0.725000 ;
      RECT 0.530000  0.725000  3.380000 0.735000 ;
      RECT 0.570000  2.175000  0.820000 2.635000 ;
      RECT 0.990000  2.005000  1.240000 2.465000 ;
      RECT 1.030000  0.085000  1.200000 0.555000 ;
      RECT 1.370000  0.255000  1.700000 0.725000 ;
      RECT 1.410000  2.175000  1.660000 2.635000 ;
      RECT 1.830000  2.005000  2.080000 2.295000 ;
      RECT 1.830000  2.295000  3.760000 2.465000 ;
      RECT 1.870000  0.085000  2.040000 0.555000 ;
      RECT 2.210000  0.255000  2.540000 0.725000 ;
      RECT 2.250000  1.615000  2.420000 1.785000 ;
      RECT 2.250000  1.785000  3.340000 1.955000 ;
      RECT 2.250000  1.955000  2.500000 2.125000 ;
      RECT 2.670000  2.125000  2.920000 2.295000 ;
      RECT 2.710000  0.085000  2.880000 0.555000 ;
      RECT 3.050000  0.255000  3.380000 0.725000 ;
      RECT 3.090000  1.955000  3.340000 2.125000 ;
      RECT 3.510000  1.795000  3.760000 2.295000 ;
      RECT 3.550000  0.085000  3.820000 0.895000 ;
      RECT 3.990000  0.255000  6.000000 0.475000 ;
      RECT 4.030000  1.785000  7.640000 2.005000 ;
      RECT 4.030000  2.005000  4.280000 2.465000 ;
      RECT 4.450000  2.175000  4.700000 2.635000 ;
      RECT 4.870000  2.005000  5.120000 2.465000 ;
      RECT 5.290000  2.175000  5.540000 2.635000 ;
      RECT 5.710000  2.005000  5.960000 2.465000 ;
      RECT 5.750000  0.475000  6.000000 0.725000 ;
      RECT 5.750000  0.725000  7.680000 0.905000 ;
      RECT 6.130000  2.175000  6.380000 2.635000 ;
      RECT 6.170000  0.085000  6.340000 0.555000 ;
      RECT 6.510000  0.255000  6.840000 0.725000 ;
      RECT 6.550000  1.455000  6.800000 1.785000 ;
      RECT 6.550000  2.005000  6.800000 2.465000 ;
      RECT 6.970000  2.175000  7.220000 2.635000 ;
      RECT 7.010000  0.085000  7.180000 0.555000 ;
      RECT 7.260000  1.445000  7.710000 1.615000 ;
      RECT 7.350000  0.255000  7.680000 0.725000 ;
      RECT 7.390000  2.005000  7.640000 2.295000 ;
      RECT 7.390000  2.295000  9.430000 2.465000 ;
      RECT 7.540000  1.105000  9.565000 1.275000 ;
      RECT 7.540000  1.275000  7.710000 1.445000 ;
      RECT 7.960000  0.085000  8.130000 0.555000 ;
      RECT 8.340000  1.835000  8.590000 2.295000 ;
      RECT 8.540000  1.075000  9.565000 1.105000 ;
      RECT 8.800000  0.085000  8.970000 0.555000 ;
      RECT 9.180000  1.795000  9.430000 2.295000 ;
      RECT 9.640000  0.085000  9.810000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  1.445000 2.155000 1.615000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  1.445000 7.675000 1.615000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 1.925000 1.415000 2.215000 1.460000 ;
      RECT 1.925000 1.460000 7.735000 1.600000 ;
      RECT 1.925000 1.600000 2.215000 1.645000 ;
      RECT 7.445000 1.415000 7.735000 1.460000 ;
      RECT 7.445000 1.600000 7.735000 1.645000 ;
  END
END sky130_fd_sc_hd__xor2_4
MACRO sky130_fd_sc_hd__or2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 0.995000 1.240000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.765000 0.345000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 0.265000 1.770000 0.735000 ;
        RECT 1.440000 0.735000 3.135000 0.905000 ;
        RECT 1.440000 1.835000 2.610000 2.005000 ;
        RECT 1.440000 2.005000 1.770000 2.465000 ;
        RECT 2.280000 0.265000 2.610000 0.735000 ;
        RECT 2.280000 1.495000 3.135000 1.665000 ;
        RECT 2.280000 1.665000 2.610000 1.835000 ;
        RECT 2.280000 2.005000 2.610000 2.465000 ;
        RECT 2.790000 0.905000 3.135000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.105000  0.085000 0.345000 0.595000 ;
      RECT 0.155000  1.495000 1.615000 1.665000 ;
      RECT 0.155000  1.665000 0.515000 2.465000 ;
      RECT 0.515000  0.290000 0.845000 0.825000 ;
      RECT 0.515000  0.825000 0.695000 1.495000 ;
      RECT 1.060000  0.085000 1.230000 0.825000 ;
      RECT 1.060000  1.835000 1.230000 2.635000 ;
      RECT 1.410000  1.075000 2.620000 1.245000 ;
      RECT 1.410000  1.245000 1.615000 1.495000 ;
      RECT 1.940000  0.085000 2.110000 0.565000 ;
      RECT 1.940000  2.175000 2.110000 2.635000 ;
      RECT 2.780000  0.085000 2.950000 0.565000 ;
      RECT 2.780000  1.835000 2.950000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__or2_4
MACRO sky130_fd_sc_hd__or2_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.995000 1.335000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.995000 0.500000 1.615000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.326800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.525000 2.180000 0.825000 ;
        RECT 1.645000 2.135000 2.180000 2.465000 ;
        RECT 1.865000 0.825000 2.180000 2.135000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.250000  0.085000 0.490000 0.825000 ;
      RECT 0.270000  1.785000 1.695000 1.955000 ;
      RECT 0.270000  1.955000 0.660000 2.130000 ;
      RECT 0.670000  0.425000 0.950000 0.825000 ;
      RECT 0.670000  0.825000 0.840000 1.785000 ;
      RECT 1.145000  2.125000 1.475000 2.635000 ;
      RECT 1.180000  0.085000 1.395000 0.825000 ;
      RECT 1.525000  0.995000 1.695000 1.785000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__or2_0
MACRO sky130_fd_sc_hd__or2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.765000 1.275000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.500000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.509000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.255000 2.180000 0.825000 ;
        RECT 1.645000 1.845000 2.180000 2.465000 ;
        RECT 1.865000 0.825000 2.180000 1.845000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.250000  0.085000 0.490000 0.595000 ;
      RECT 0.270000  1.495000 1.695000 1.665000 ;
      RECT 0.270000  1.665000 0.660000 1.840000 ;
      RECT 0.670000  0.265000 0.950000 0.595000 ;
      RECT 0.670000  0.595000 0.840000 1.495000 ;
      RECT 1.145000  1.835000 1.475000 2.635000 ;
      RECT 1.180000  0.085000 1.395000 0.595000 ;
      RECT 1.525000  0.995000 1.695000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__or2_1
MACRO sky130_fd_sc_hd__or2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 0.765000 1.275000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.765000 0.345000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.440000 1.835000 2.215000 2.005000 ;
        RECT 1.440000 2.005000 1.770000 2.465000 ;
        RECT 1.520000 0.385000 1.690000 0.655000 ;
        RECT 1.520000 0.655000 2.215000 0.825000 ;
        RECT 1.785000 0.825000 2.215000 1.835000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.105000  0.085000 0.345000 0.595000 ;
      RECT 0.155000  1.495000 1.615000 1.665000 ;
      RECT 0.155000  1.665000 0.515000 1.840000 ;
      RECT 0.515000  0.255000 0.805000 0.595000 ;
      RECT 0.515000  0.595000 0.695000 1.495000 ;
      RECT 1.035000  0.085000 1.350000 0.595000 ;
      RECT 1.100000  1.835000 1.270000 2.635000 ;
      RECT 1.445000  0.995000 1.615000 1.495000 ;
      RECT 1.860000  0.085000 2.190000 0.485000 ;
      RECT 1.940000  2.175000 2.110000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__or2_2
MACRO sky130_fd_sc_hd__clkdlybuf4s25_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s25_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.495000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.497000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.770000 0.285000 3.095000 0.615000 ;
        RECT 2.770000 1.625000 3.095000 2.460000 ;
        RECT 2.865000 0.615000 3.095000 0.765000 ;
        RECT 2.865000 0.765000 3.595000 1.275000 ;
        RECT 2.865000 1.275000 3.095000 1.625000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  0.305000 0.345000 0.640000 ;
      RECT 0.095000  0.640000 0.840000 0.810000 ;
      RECT 0.095000  1.785000 0.835000 1.955000 ;
      RECT 0.095000  1.955000 0.345000 2.465000 ;
      RECT 0.575000  0.085000 0.905000 0.470000 ;
      RECT 0.575000  2.125000 0.905000 2.635000 ;
      RECT 0.665000  0.810000 0.840000 0.995000 ;
      RECT 0.665000  0.995000 1.035000 1.325000 ;
      RECT 0.665000  1.325000 1.005000 1.750000 ;
      RECT 0.665000  1.750000 0.835000 1.785000 ;
      RECT 1.095000  0.255000 1.425000 0.780000 ;
      RECT 1.175000  1.425000 1.440000 2.465000 ;
      RECT 1.205000  0.780000 1.425000 0.995000 ;
      RECT 1.205000  0.995000 2.165000 1.325000 ;
      RECT 1.205000  1.325000 1.440000 1.425000 ;
      RECT 1.615000  0.255000 1.945000 0.635000 ;
      RECT 1.615000  0.635000 2.595000 0.805000 ;
      RECT 1.695000  1.500000 2.595000 1.745000 ;
      RECT 1.695000  1.745000 1.945000 2.465000 ;
      RECT 2.135000  0.085000 2.465000 0.465000 ;
      RECT 2.135000  1.915000 2.465000 2.635000 ;
      RECT 2.335000  0.805000 2.595000 1.500000 ;
      RECT 3.265000  0.085000 3.595000 0.550000 ;
      RECT 3.265000  1.635000 3.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s25_2
MACRO sky130_fd_sc_hd__clkdlybuf4s25_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s25_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.485000 1.320000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.702900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.015000 0.255000 3.595000 0.640000 ;
        RECT 3.035000 1.565000 3.595000 2.465000 ;
        RECT 3.230000 0.640000 3.595000 1.565000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.255000 0.410000 0.735000 ;
      RECT 0.085000  0.735000 1.005000 0.905000 ;
      RECT 0.085000  1.490000 1.005000 1.660000 ;
      RECT 0.085000  1.660000 0.430000 2.465000 ;
      RECT 0.580000  0.085000 0.910000 0.565000 ;
      RECT 0.600000  1.830000 0.925000 2.635000 ;
      RECT 0.655000  0.905000 1.005000 1.025000 ;
      RECT 0.655000  1.025000 1.105000 1.295000 ;
      RECT 0.655000  1.295000 1.005000 1.490000 ;
      RECT 1.175000  0.255000 1.645000 0.855000 ;
      RECT 1.195000  1.790000 1.645000 2.465000 ;
      RECT 1.470000  0.855000 1.645000 1.075000 ;
      RECT 1.470000  1.075000 2.420000 1.250000 ;
      RECT 1.470000  1.250000 1.645000 1.790000 ;
      RECT 1.815000  0.255000 2.065000 0.735000 ;
      RECT 1.815000  0.735000 2.765000 0.905000 ;
      RECT 1.815000  1.495000 2.765000 1.665000 ;
      RECT 1.815000  1.665000 2.065000 2.465000 ;
      RECT 2.235000  1.835000 2.845000 2.635000 ;
      RECT 2.240000  0.085000 2.845000 0.565000 ;
      RECT 2.595000  0.905000 2.765000 0.990000 ;
      RECT 2.595000  0.990000 3.050000 1.325000 ;
      RECT 2.595000  1.325000 2.765000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s25_1
MACRO sky130_fd_sc_hd__nand4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 1.075000 4.495000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.235000 1.075000 3.080000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.075000 1.700000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.845000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.445000 3.925000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 2.355000 1.665000 2.685000 2.465000 ;
        RECT 3.370000 1.055000 3.925000 1.445000 ;
        RECT 3.595000 0.635000 3.925000 1.055000 ;
        RECT 3.595000 1.665000 3.925000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 1.185000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 0.935000  0.255000 2.125000 0.465000 ;
      RECT 0.935000  0.465000 1.185000 0.735000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.355000  0.635000 3.085000 0.905000 ;
      RECT 1.855000  1.835000 2.185000 2.635000 ;
      RECT 2.315000  0.255000 4.425000 0.465000 ;
      RECT 2.995000  1.835000 3.325000 2.635000 ;
      RECT 3.255000  0.465000 3.425000 0.885000 ;
      RECT 4.095000  0.465000 4.425000 0.905000 ;
      RECT 4.095000  1.445000 4.425000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4_2
MACRO sky130_fd_sc_hd__nand4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 0.995000 2.215000 1.665000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.300000 1.350000 0.825000 ;
        RECT 1.145000 0.825000 1.350000 0.995000 ;
        RECT 1.145000 0.995000 1.455000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.300000 0.810000 0.995000 ;
        RECT 0.595000 0.995000 0.975000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.995000 0.395000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.795000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.495000 1.795000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.385000 1.665000 1.715000 2.465000 ;
        RECT 1.520000 0.255000 2.215000 0.825000 ;
        RECT 1.625000 0.825000 1.795000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.090000  0.085000 0.425000 0.825000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4_1
MACRO sky130_fd_sc_hd__nand4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465000 1.075000 7.710000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.850000 1.075000 5.565000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.075000 3.540000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.700000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.445000 7.305000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 2.195000 1.665000 2.525000 2.465000 ;
        RECT 3.035000 1.665000 3.365000 2.465000 ;
        RECT 4.395000 1.665000 4.725000 2.465000 ;
        RECT 5.235000 1.665000 5.565000 2.465000 ;
        RECT 6.110000 0.655000 7.305000 0.905000 ;
        RECT 6.110000 0.905000 6.290000 1.445000 ;
        RECT 6.135000 1.665000 6.465000 2.465000 ;
        RECT 6.975000 1.665000 7.305000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.090000  0.255000 0.345000 0.655000 ;
      RECT 0.090000  0.655000 2.025000 0.905000 ;
      RECT 0.090000  1.445000 0.345000 2.635000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 1.015000  0.255000 1.185000 0.655000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.355000  0.085000 1.685000 0.485000 ;
      RECT 1.855000  0.255000 3.785000 0.485000 ;
      RECT 1.855000  0.485000 2.025000 0.655000 ;
      RECT 1.855000  1.835000 2.025000 2.635000 ;
      RECT 2.195000  0.655000 5.565000 0.905000 ;
      RECT 2.695000  1.835000 2.865000 2.635000 ;
      RECT 3.535000  1.835000 4.225000 2.635000 ;
      RECT 3.975000  0.255000 7.730000 0.485000 ;
      RECT 4.895000  1.835000 5.065000 2.635000 ;
      RECT 5.770000  0.485000 5.940000 0.905000 ;
      RECT 5.770000  1.835000 5.940000 2.635000 ;
      RECT 6.635000  1.835000 6.805000 2.635000 ;
      RECT 7.475000  0.485000 7.730000 0.905000 ;
      RECT 7.475000  1.445000 7.735000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4_4
MACRO sky130_fd_sc_hd__ha_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ha_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 1.055000 4.045000 1.225000 ;
        RECT 3.820000 1.225000 4.045000 1.675000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.310000 1.005000 2.615000 1.395000 ;
        RECT 2.310000 1.395000 3.595000 1.675000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635000 0.315000 4.965000 0.825000 ;
        RECT 4.715000 1.545000 4.965000 2.415000 ;
        RECT 4.790000 0.825000 4.965000 1.545000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.315000 0.885000 0.825000 ;
        RECT 0.555000 0.825000 0.780000 1.565000 ;
        RECT 0.555000 1.565000 0.885000 2.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.135000  0.085000 0.375000 0.885000 ;
      RECT 0.135000  1.495000 0.375000 2.635000 ;
      RECT 0.950000  1.075000 1.590000 1.245000 ;
      RECT 1.055000  0.085000 1.250000 0.885000 ;
      RECT 1.055000  1.515000 1.250000 2.635000 ;
      RECT 1.420000  0.345000 1.745000 0.675000 ;
      RECT 1.420000  0.675000 1.590000 1.075000 ;
      RECT 1.420000  1.245000 1.590000 2.205000 ;
      RECT 1.420000  2.205000 2.220000 2.375000 ;
      RECT 1.760000  0.995000 1.930000 1.855000 ;
      RECT 1.760000  1.855000 4.465000 2.025000 ;
      RECT 1.995000  0.345000 2.165000 0.635000 ;
      RECT 1.995000  0.635000 3.005000 0.805000 ;
      RECT 2.335000  0.085000 2.665000 0.465000 ;
      RECT 2.835000  0.345000 3.005000 0.635000 ;
      RECT 2.850000  2.205000 3.640000 2.635000 ;
      RECT 3.460000  0.345000 3.630000 0.715000 ;
      RECT 3.460000  0.715000 4.465000 0.885000 ;
      RECT 3.810000  2.025000 3.980000 2.355000 ;
      RECT 4.215000  0.085000 4.465000 0.545000 ;
      RECT 4.215000  2.205000 4.545000 2.635000 ;
      RECT 4.295000  0.885000 4.465000 0.995000 ;
      RECT 4.295000  0.995000 4.620000 1.325000 ;
      RECT 4.295000  1.325000 4.465000 1.855000 ;
      RECT 5.145000  0.085000 5.385000 0.885000 ;
      RECT 5.145000  1.495000 5.385000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__ha_2
MACRO sky130_fd_sc_hd__ha_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ha_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335000 1.315000 3.585000 1.485000 ;
        RECT 3.360000 1.055000 3.585000 1.315000 ;
        RECT 3.360000 1.485000 3.585000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.850000 1.345000 2.155000 1.655000 ;
        RECT 1.850000 1.655000 3.165000 1.825000 ;
        RECT 1.850000 1.825000 2.155000 2.375000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 0.315000 4.515000 0.825000 ;
        RECT 4.175000 1.565000 4.515000 2.415000 ;
        RECT 4.330000 0.825000 4.515000 1.565000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.315000 0.425000 0.825000 ;
        RECT 0.090000 0.825000 0.320000 1.565000 ;
        RECT 0.090000 1.565000 0.425000 2.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.490000  1.075000 1.130000 1.245000 ;
      RECT 0.595000  0.085000 0.790000 0.885000 ;
      RECT 0.595000  1.515000 0.790000 2.275000 ;
      RECT 0.595000  2.275000 1.260000 2.635000 ;
      RECT 0.960000  0.345000 1.285000 0.675000 ;
      RECT 0.960000  0.675000 1.130000 1.075000 ;
      RECT 0.960000  1.245000 1.130000 1.935000 ;
      RECT 0.960000  1.935000 1.680000 2.105000 ;
      RECT 1.300000  0.975000 3.170000 1.145000 ;
      RECT 1.300000  1.145000 1.470000 1.325000 ;
      RECT 1.510000  2.105000 1.680000 2.355000 ;
      RECT 1.535000  0.345000 1.705000 0.635000 ;
      RECT 1.535000  0.635000 2.545000 0.805000 ;
      RECT 1.875000  0.085000 2.205000 0.465000 ;
      RECT 2.375000  0.345000 2.545000 0.635000 ;
      RECT 2.450000  2.275000 3.120000 2.635000 ;
      RECT 3.000000  0.345000 3.170000 0.715000 ;
      RECT 3.000000  0.715000 4.005000 0.885000 ;
      RECT 3.000000  0.885000 3.170000 0.975000 ;
      RECT 3.350000  1.785000 4.005000 1.955000 ;
      RECT 3.350000  1.955000 3.520000 2.355000 ;
      RECT 3.755000  0.085000 4.005000 0.545000 ;
      RECT 3.755000  2.125000 4.005000 2.635000 ;
      RECT 3.835000  0.885000 4.005000 0.995000 ;
      RECT 3.835000  0.995000 4.160000 1.325000 ;
      RECT 3.835000  1.325000 4.005000 1.785000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__ha_1
MACRO sky130_fd_sc_hd__ha_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ha_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.320000 1.075000 4.380000 1.245000 ;
        RECT 4.210000 1.245000 4.380000 1.505000 ;
        RECT 4.210000 1.505000 6.810000 1.675000 ;
        RECT 5.625000 0.995000 5.795000 1.505000 ;
        RECT 6.580000 0.995000 7.055000 1.325000 ;
        RECT 6.580000 1.325000 6.810000 1.505000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.550000 0.995000 5.455000 1.165000 ;
        RECT 4.550000 1.165000 4.720000 1.325000 ;
        RECT 5.285000 0.730000 6.315000 0.825000 ;
        RECT 5.285000 0.825000 5.535000 0.845000 ;
        RECT 5.285000 0.845000 5.495000 0.875000 ;
        RECT 5.285000 0.875000 5.455000 0.995000 ;
        RECT 5.295000 0.720000 6.315000 0.730000 ;
        RECT 5.310000 0.710000 6.315000 0.720000 ;
        RECT 5.320000 0.695000 6.315000 0.710000 ;
        RECT 5.335000 0.675000 6.315000 0.695000 ;
        RECT 5.345000 0.655000 6.315000 0.675000 ;
        RECT 6.085000 0.825000 6.315000 1.325000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.595000 0.315000 7.845000 0.735000 ;
        RECT 7.595000 0.735000 8.685000 0.905000 ;
        RECT 7.595000 1.415000 8.685000 1.585000 ;
        RECT 7.595000 1.585000 7.765000 2.415000 ;
        RECT 8.405000 0.315000 8.685000 0.735000 ;
        RECT 8.405000 0.905000 8.685000 1.415000 ;
        RECT 8.405000 1.585000 8.685000 2.415000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.315000 0.845000 1.065000 ;
        RECT 0.515000 1.065000 1.550000 1.335000 ;
        RECT 0.515000 1.335000 0.845000 2.415000 ;
        RECT 1.355000 0.315000 1.685000 0.825000 ;
        RECT 1.355000 0.825000 1.550000 1.065000 ;
        RECT 1.355000 1.335000 1.550000 1.565000 ;
        RECT 1.355000 1.565000 1.685000 2.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.135000  0.085000 0.345000 0.885000 ;
      RECT 0.135000  1.495000 0.345000 2.635000 ;
      RECT 1.015000  0.085000 1.185000 0.885000 ;
      RECT 1.015000  1.515000 1.185000 2.635000 ;
      RECT 1.720000  1.075000 2.750000 1.245000 ;
      RECT 1.855000  0.085000 2.095000 0.885000 ;
      RECT 1.855000  1.495000 2.365000 2.635000 ;
      RECT 2.270000  0.305000 3.385000 0.475000 ;
      RECT 2.580000  0.645000 3.045000 0.815000 ;
      RECT 2.580000  0.815000 2.750000 1.075000 ;
      RECT 2.580000  1.245000 2.750000 1.765000 ;
      RECT 2.580000  1.765000 3.700000 1.935000 ;
      RECT 2.770000  1.935000 2.940000 2.355000 ;
      RECT 2.920000  0.995000 3.090000 1.425000 ;
      RECT 2.920000  1.425000 4.040000 1.595000 ;
      RECT 3.190000  2.105000 3.360000 2.635000 ;
      RECT 3.215000  0.475000 3.385000 0.645000 ;
      RECT 3.215000  0.645000 5.115000 0.815000 ;
      RECT 3.530000  1.935000 3.700000 2.205000 ;
      RECT 3.530000  2.205000 4.330000 2.375000 ;
      RECT 3.555000  0.085000 3.910000 0.465000 ;
      RECT 3.870000  1.595000 4.040000 1.855000 ;
      RECT 3.870000  1.855000 7.395000 2.025000 ;
      RECT 4.080000  0.345000 4.250000 0.645000 ;
      RECT 4.420000  0.085000 4.750000 0.465000 ;
      RECT 4.920000  0.255000 5.190000 0.585000 ;
      RECT 4.920000  0.585000 5.115000 0.645000 ;
      RECT 5.240000  2.205000 5.570000 2.635000 ;
      RECT 5.385000  0.085000 5.715000 0.465000 ;
      RECT 5.835000  2.025000 6.005000 2.355000 ;
      RECT 6.175000  0.295000 6.875000 0.465000 ;
      RECT 6.175000  2.205000 6.505000 2.635000 ;
      RECT 6.675000  2.025000 6.845000 2.355000 ;
      RECT 6.705000  0.465000 6.875000 0.645000 ;
      RECT 6.705000  0.645000 7.395000 0.815000 ;
      RECT 7.055000  0.085000 7.385000 0.465000 ;
      RECT 7.055000  2.205000 7.385000 2.635000 ;
      RECT 7.225000  0.815000 7.395000 1.075000 ;
      RECT 7.225000  1.075000 8.225000 1.245000 ;
      RECT 7.225000  1.245000 7.395000 1.855000 ;
      RECT 7.935000  1.755000 8.225000 2.635000 ;
      RECT 8.015000  0.085000 8.225000 0.565000 ;
      RECT 8.855000  0.085000 9.065000 0.885000 ;
      RECT 8.855000  1.495000 9.065000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
END sky130_fd_sc_hd__ha_4
MACRO sky130_fd_sc_hd__nand4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.995000 0.330000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 0.995000 0.975000 1.615000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.120000 1.075000 7.910000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.420000 1.075000 10.015000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.540000 0.655000 3.990000 0.905000 ;
        RECT 2.540000 1.445000 9.590000 1.665000 ;
        RECT 2.540000 1.665000 2.790000 2.465000 ;
        RECT 3.380000 1.665000 3.710000 2.465000 ;
        RECT 3.700000 0.905000 3.990000 1.445000 ;
        RECT 4.220000 1.665000 4.550000 2.465000 ;
        RECT 5.060000 1.665000 5.390000 2.465000 ;
        RECT 6.740000 1.665000 7.070000 2.465000 ;
        RECT 7.580000 1.665000 7.910000 2.465000 ;
        RECT 8.420000 1.665000 8.750000 2.465000 ;
        RECT 9.260000 1.665000 9.590000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.255000  0.345000 0.635000 ;
      RECT 0.085000  0.635000  1.455000 0.805000 ;
      RECT 0.085000  1.785000  1.455000 1.980000 ;
      RECT 0.085000  1.980000  0.370000 2.440000 ;
      RECT 0.515000  0.085000  0.845000 0.465000 ;
      RECT 0.540000  2.195000  0.765000 2.635000 ;
      RECT 0.935000  2.150000  1.795000 2.465000 ;
      RECT 1.015000  0.255000  1.795000 0.465000 ;
      RECT 1.145000  0.805000  1.455000 1.785000 ;
      RECT 1.625000  0.465000  1.795000 1.075000 ;
      RECT 1.625000  1.075000  2.210000 1.305000 ;
      RECT 1.625000  1.305000  1.795000 2.150000 ;
      RECT 2.200000  0.255000  5.810000 0.485000 ;
      RECT 2.200000  0.485000  2.370000 0.905000 ;
      RECT 2.200000  1.495000  2.370000 2.635000 ;
      RECT 2.540000  1.075000  3.285000 1.245000 ;
      RECT 2.960000  1.835000  3.210000 2.635000 ;
      RECT 3.880000  1.835000  4.050000 2.635000 ;
      RECT 4.160000  1.075000  5.390000 1.275000 ;
      RECT 4.220000  0.655000  5.390000 0.735000 ;
      RECT 4.220000  0.735000  6.150000 0.905000 ;
      RECT 4.720000  1.835000  4.890000 2.635000 ;
      RECT 5.610000  1.835000  6.540000 2.635000 ;
      RECT 5.980000  0.255000  7.910000 0.485000 ;
      RECT 5.980000  0.485000  6.150000 0.735000 ;
      RECT 6.320000  0.655000 10.035000 0.905000 ;
      RECT 7.240000  1.835000  7.410000 2.635000 ;
      RECT 8.080000  1.835000  8.250000 2.635000 ;
      RECT 8.420000  0.085000  8.750000 0.485000 ;
      RECT 8.920000  1.835000  9.090000 2.635000 ;
      RECT 9.260000  0.085000  9.590000 0.485000 ;
      RECT 9.760000  1.445000 10.035000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.980000  1.105000 2.150000 1.275000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.280000  1.105000 4.450000 1.275000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 1.920000 1.075000 2.210000 1.120000 ;
      RECT 1.920000 1.120000 4.510000 1.260000 ;
      RECT 1.920000 1.260000 2.210000 1.305000 ;
      RECT 4.220000 1.075000 4.510000 1.120000 ;
      RECT 4.220000 1.260000 4.510000 1.305000 ;
  END
END sky130_fd_sc_hd__nand4bb_4
MACRO sky130_fd_sc_hd__nand4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.390000 0.725000 3.640000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.075000 0.780000 1.655000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 0.735000 1.720000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.970000 1.075000 1.320000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.909000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.120000 1.495000 2.670000 1.665000 ;
        RECT 1.120000 1.665000 1.450000 2.465000 ;
        RECT 2.140000 1.665000 2.470000 2.465000 ;
        RECT 2.420000 0.255000 2.930000 0.825000 ;
        RECT 2.420000 0.825000 2.670000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.485000 0.425000 0.715000 ;
      RECT 0.085000  0.715000 1.270000 0.905000 ;
      RECT 0.085000  0.905000 0.260000 2.065000 ;
      RECT 0.085000  2.065000 0.425000 2.465000 ;
      RECT 0.595000  0.085000 0.900000 0.545000 ;
      RECT 0.595000  1.835000 0.925000 2.635000 ;
      RECT 1.080000  0.365000 2.250000 0.555000 ;
      RECT 1.080000  0.555000 1.270000 0.715000 ;
      RECT 1.640000  1.835000 1.970000 2.635000 ;
      RECT 1.970000  0.555000 2.250000 1.325000 ;
      RECT 2.680000  2.175000 3.450000 2.635000 ;
      RECT 2.840000  0.995000 3.090000 1.835000 ;
      RECT 2.840000  1.835000 4.055000 2.005000 ;
      RECT 3.100000  0.085000 3.450000 0.545000 ;
      RECT 3.620000  0.255000 4.055000 0.545000 ;
      RECT 3.635000  2.005000 4.055000 2.465000 ;
      RECT 3.810000  0.545000 4.055000 1.835000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__nand4bb_1
MACRO sky130_fd_sc_hd__nand4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.170000 0.890000 1.340000 ;
        RECT 0.610000 1.070000 0.890000 1.170000 ;
        RECT 0.610000 1.340000 0.890000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.070000 0.330000 1.615000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.720000 1.075000 4.615000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.945000 1.075000 5.875000 1.275000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.085000 0.655000 2.415000 1.445000 ;
        RECT 2.085000 1.445000 5.455000 1.665000 ;
        RECT 2.085000 1.665000 2.335000 2.465000 ;
        RECT 2.925000 1.665000 3.255000 2.465000 ;
        RECT 3.245000 1.075000 3.550000 1.445000 ;
        RECT 4.285000 1.665000 4.615000 2.465000 ;
        RECT 5.125000 1.665000 5.455000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.730000 ;
      RECT 0.085000  0.730000 1.230000 0.900000 ;
      RECT 0.085000  1.785000 1.230000 1.980000 ;
      RECT 0.085000  1.980000 0.370000 2.440000 ;
      RECT 0.515000  0.085000 0.765000 0.545000 ;
      RECT 0.540000  2.195000 0.765000 2.635000 ;
      RECT 0.935000  0.255000 1.575000 0.560000 ;
      RECT 0.935000  2.150000 1.575000 2.465000 ;
      RECT 1.060000  0.900000 1.230000 1.785000 ;
      RECT 1.400000  0.560000 1.575000 0.715000 ;
      RECT 1.400000  0.715000 1.580000 1.410000 ;
      RECT 1.400000  1.410000 1.575000 2.150000 ;
      RECT 1.745000  0.255000 3.675000 0.485000 ;
      RECT 1.745000  0.485000 1.915000 0.585000 ;
      RECT 1.745000  1.495000 1.915000 2.635000 ;
      RECT 2.505000  1.835000 2.755000 2.635000 ;
      RECT 2.745000  1.075000 3.075000 1.275000 ;
      RECT 2.925000  0.655000 4.615000 0.905000 ;
      RECT 3.425000  1.835000 4.115000 2.635000 ;
      RECT 3.865000  0.255000 5.035000 0.485000 ;
      RECT 4.785000  0.485000 5.035000 0.735000 ;
      RECT 4.785000  0.735000 5.895000 0.905000 ;
      RECT 4.785000  1.835000 4.955000 2.635000 ;
      RECT 5.205000  0.085000 5.375000 0.565000 ;
      RECT 5.545000  0.255000 5.895000 0.735000 ;
      RECT 5.625000  1.445000 5.895000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.060000  1.105000 1.230000 1.275000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  1.105000 3.075000 1.275000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 1.000000 1.075000 3.135000 1.305000 ;
  END
END sky130_fd_sc_hd__nand4bb_2
MACRO sky130_fd_sc_hd__dfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfsbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.005000 2.180000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.865000 0.255000 10.125000 0.825000 ;
        RECT 9.865000 1.445000 10.125000 2.465000 ;
        RECT 9.910000 0.825000 10.125000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.370000 0.255000 8.700000 2.465000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 0.735000 4.020000 1.065000 ;
      LAYER mcon ;
        RECT 3.825000 0.765000 3.995000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.660000 0.735000 7.320000 1.005000 ;
        RECT 6.660000 1.005000 6.990000 1.065000 ;
      LAYER mcon ;
        RECT 7.045000 0.765000 7.215000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765000 0.735000 4.055000 0.780000 ;
        RECT 3.765000 0.780000 7.275000 0.920000 ;
        RECT 3.765000 0.920000 4.055000 0.965000 ;
        RECT 6.985000 0.735000 7.275000 0.780000 ;
        RECT 6.985000 0.920000 7.275000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.770000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.580000 0.085000 ;
      RECT 0.000000  2.635000 10.580000 2.805000 ;
      RECT 0.175000  0.345000  0.345000 0.635000 ;
      RECT 0.175000  0.635000  0.840000 0.805000 ;
      RECT 0.175000  1.795000  0.840000 1.965000 ;
      RECT 0.175000  1.965000  0.345000 2.465000 ;
      RECT 0.515000  0.085000  0.845000 0.465000 ;
      RECT 0.515000  2.135000  0.845000 2.635000 ;
      RECT 0.610000  0.805000  0.840000 1.795000 ;
      RECT 1.015000  0.345000  1.240000 2.465000 ;
      RECT 1.430000  0.635000  2.125000 0.825000 ;
      RECT 1.430000  0.825000  1.600000 1.795000 ;
      RECT 1.430000  1.795000  2.125000 1.965000 ;
      RECT 1.455000  0.085000  1.785000 0.465000 ;
      RECT 1.455000  2.135000  1.785000 2.635000 ;
      RECT 1.955000  0.305000  2.125000 0.635000 ;
      RECT 1.955000  1.965000  2.125000 2.465000 ;
      RECT 2.350000  0.705000  2.570000 1.575000 ;
      RECT 2.350000  1.575000  2.850000 1.955000 ;
      RECT 2.360000  2.250000  3.190000 2.420000 ;
      RECT 2.425000  0.265000  3.440000 0.465000 ;
      RECT 2.750000  0.645000  3.100000 1.015000 ;
      RECT 3.020000  1.195000  3.440000 1.235000 ;
      RECT 3.020000  1.235000  4.370000 1.405000 ;
      RECT 3.020000  1.405000  3.190000 2.250000 ;
      RECT 3.270000  0.465000  3.440000 1.195000 ;
      RECT 3.360000  1.575000  3.610000 1.835000 ;
      RECT 3.360000  1.835000  4.710000 2.085000 ;
      RECT 3.430000  2.255000  3.810000 2.635000 ;
      RECT 3.610000  0.085000  4.020000 0.525000 ;
      RECT 3.990000  2.085000  4.160000 2.375000 ;
      RECT 4.120000  1.405000  4.370000 1.565000 ;
      RECT 4.310000  0.295000  4.560000 0.725000 ;
      RECT 4.310000  0.725000  4.710000 1.065000 ;
      RECT 4.330000  2.255000  4.660000 2.635000 ;
      RECT 4.540000  1.065000  4.710000 1.835000 ;
      RECT 4.740000  0.085000  5.080000 0.545000 ;
      RECT 4.900000  0.725000  6.150000 0.895000 ;
      RECT 4.900000  0.895000  5.070000 1.655000 ;
      RECT 4.900000  1.655000  5.400000 1.965000 ;
      RECT 5.110000  2.165000  5.760000 2.415000 ;
      RECT 5.240000  1.065000  5.420000 1.475000 ;
      RECT 5.590000  1.235000  7.470000 1.405000 ;
      RECT 5.590000  1.405000  5.760000 1.915000 ;
      RECT 5.590000  1.915000  6.780000 2.085000 ;
      RECT 5.590000  2.085000  5.760000 2.165000 ;
      RECT 5.640000  0.305000  6.490000 0.475000 ;
      RECT 5.820000  0.895000  6.150000 1.015000 ;
      RECT 5.930000  1.575000  7.830000 1.745000 ;
      RECT 5.930000  2.255000  6.340000 2.635000 ;
      RECT 6.320000  0.475000  6.490000 1.235000 ;
      RECT 6.540000  2.085000  6.780000 2.375000 ;
      RECT 6.670000  0.085000  7.330000 0.565000 ;
      RECT 7.010000  1.945000  7.340000 2.635000 ;
      RECT 7.140000  1.175000  7.470000 1.235000 ;
      RECT 7.510000  0.350000  7.830000 0.680000 ;
      RECT 7.510000  1.745000  7.830000 1.765000 ;
      RECT 7.510000  1.765000  7.680000 2.375000 ;
      RECT 7.640000  0.680000  7.830000 1.575000 ;
      RECT 8.020000  0.085000  8.200000 0.905000 ;
      RECT 8.020000  1.480000  8.200000 2.635000 ;
      RECT 8.890000  0.255000  9.220000 0.995000 ;
      RECT 8.890000  0.995000  9.740000 1.325000 ;
      RECT 8.890000  1.325000  9.220000 2.465000 ;
      RECT 9.445000  0.085000  9.615000 0.585000 ;
      RECT 9.445000  1.825000  9.615000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.645000  1.785000  0.815000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  0.765000  1.235000 0.935000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.785000  2.615000 1.955000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  0.765000  3.075000 0.935000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.245000  1.105000  5.415000 1.275000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 5.435000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 1.005000 0.735000 1.295000 0.780000 ;
      RECT 1.005000 0.780000 3.135000 0.920000 ;
      RECT 1.005000 0.920000 1.295000 0.965000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.845000 0.735000 3.135000 0.780000 ;
      RECT 2.845000 0.920000 3.135000 0.965000 ;
      RECT 2.920000 0.965000 3.135000 1.120000 ;
      RECT 2.920000 1.120000 5.475000 1.260000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 5.185000 1.075000 5.475000 1.120000 ;
      RECT 5.185000 1.260000 5.475000 1.305000 ;
  END
END sky130_fd_sc_hd__dfsbp_1
MACRO sky130_fd_sc_hd__dfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfsbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.005000 2.180000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.150000 1.495000 10.915000 1.665000 ;
        RECT 10.150000 1.665000 10.480000 2.465000 ;
        RECT 10.230000 0.255000 10.480000 0.720000 ;
        RECT 10.230000 0.720000 10.915000 0.825000 ;
        RECT 10.345000 0.825000 10.915000 0.845000 ;
        RECT 10.360000 0.845000 10.915000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.370000 0.255000 8.700000 2.465000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 0.735000 4.020000 1.065000 ;
      LAYER mcon ;
        RECT 3.825000 0.765000 3.995000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.660000 0.735000 7.320000 1.005000 ;
        RECT 6.660000 1.005000 6.990000 1.065000 ;
      LAYER mcon ;
        RECT 7.045000 0.765000 7.215000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765000 0.735000 4.055000 0.780000 ;
        RECT 3.765000 0.780000 7.275000 0.920000 ;
        RECT 3.765000 0.920000 4.055000 0.965000 ;
        RECT 6.985000 0.735000 7.275000 0.780000 ;
        RECT 6.985000 0.920000 7.275000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.840000 0.805000 ;
      RECT  0.175000  1.795000  0.840000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.240000 2.465000 ;
      RECT  1.430000  0.635000  2.125000 0.825000 ;
      RECT  1.430000  0.825000  1.600000 1.795000 ;
      RECT  1.430000  1.795000  2.125000 1.965000 ;
      RECT  1.455000  0.085000  1.785000 0.465000 ;
      RECT  1.455000  2.135000  1.785000 2.635000 ;
      RECT  1.955000  0.305000  2.125000 0.635000 ;
      RECT  1.955000  1.965000  2.125000 2.465000 ;
      RECT  2.350000  0.705000  2.570000 1.575000 ;
      RECT  2.350000  1.575000  2.850000 1.955000 ;
      RECT  2.360000  2.250000  3.190000 2.420000 ;
      RECT  2.425000  0.265000  3.440000 0.465000 ;
      RECT  2.750000  0.645000  3.100000 1.015000 ;
      RECT  3.020000  1.195000  3.440000 1.235000 ;
      RECT  3.020000  1.235000  4.370000 1.405000 ;
      RECT  3.020000  1.405000  3.190000 2.250000 ;
      RECT  3.270000  0.465000  3.440000 1.195000 ;
      RECT  3.360000  1.575000  3.610000 1.835000 ;
      RECT  3.360000  1.835000  4.710000 2.085000 ;
      RECT  3.430000  2.255000  3.810000 2.635000 ;
      RECT  3.610000  0.085000  4.020000 0.525000 ;
      RECT  3.990000  2.085000  4.160000 2.375000 ;
      RECT  4.120000  1.405000  4.370000 1.565000 ;
      RECT  4.310000  0.295000  4.560000 0.725000 ;
      RECT  4.310000  0.725000  4.710000 1.065000 ;
      RECT  4.330000  2.255000  4.660000 2.635000 ;
      RECT  4.540000  1.065000  4.710000 1.835000 ;
      RECT  4.740000  0.085000  5.080000 0.545000 ;
      RECT  4.900000  0.725000  6.150000 0.895000 ;
      RECT  4.900000  0.895000  5.070000 1.655000 ;
      RECT  4.900000  1.655000  5.400000 1.965000 ;
      RECT  5.110000  2.165000  5.760000 2.415000 ;
      RECT  5.240000  1.065000  5.420000 1.475000 ;
      RECT  5.590000  1.235000  7.470000 1.405000 ;
      RECT  5.590000  1.405000  5.760000 1.915000 ;
      RECT  5.590000  1.915000  6.780000 2.085000 ;
      RECT  5.590000  2.085000  5.760000 2.165000 ;
      RECT  5.640000  0.305000  6.490000 0.475000 ;
      RECT  5.820000  0.895000  6.150000 1.015000 ;
      RECT  5.930000  1.575000  7.830000 1.745000 ;
      RECT  5.930000  2.255000  6.340000 2.635000 ;
      RECT  6.320000  0.475000  6.490000 1.235000 ;
      RECT  6.540000  2.085000  6.780000 2.375000 ;
      RECT  6.670000  0.085000  7.330000 0.565000 ;
      RECT  7.010000  1.945000  7.340000 2.635000 ;
      RECT  7.140000  1.175000  7.470000 1.235000 ;
      RECT  7.510000  0.350000  7.830000 0.680000 ;
      RECT  7.510000  1.745000  7.830000 1.765000 ;
      RECT  7.510000  1.765000  7.680000 2.375000 ;
      RECT  7.640000  0.680000  7.830000 1.575000 ;
      RECT  8.020000  0.085000  8.200000 0.905000 ;
      RECT  8.020000  1.480000  8.200000 2.635000 ;
      RECT  8.870000  0.085000  9.120000 0.905000 ;
      RECT  8.870000  1.480000  9.120000 2.635000 ;
      RECT  9.310000  0.255000  9.560000 0.995000 ;
      RECT  9.310000  0.995000 10.190000 1.325000 ;
      RECT  9.310000  1.325000  9.640000 2.465000 ;
      RECT  9.730000  0.085000 10.060000 0.825000 ;
      RECT  9.810000  1.495000  9.980000 2.635000 ;
      RECT 10.650000  0.085000 10.915000 0.550000 ;
      RECT 10.650000  1.835000 10.915000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.645000  1.785000  0.815000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  0.765000  1.235000 0.935000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.785000  2.615000 1.955000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  0.765000  3.075000 0.935000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.245000  1.105000  5.415000 1.275000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 5.435000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 1.005000 0.735000 1.295000 0.780000 ;
      RECT 1.005000 0.780000 3.135000 0.920000 ;
      RECT 1.005000 0.920000 1.295000 0.965000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.845000 0.735000 3.135000 0.780000 ;
      RECT 2.845000 0.920000 3.135000 0.965000 ;
      RECT 2.920000 0.965000 3.135000 1.120000 ;
      RECT 2.920000 1.120000 5.475000 1.260000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 5.185000 1.075000 5.475000 1.120000 ;
      RECT 5.185000 1.260000 5.475000 1.305000 ;
  END
END sky130_fd_sc_hd__dfsbp_2
MACRO sky130_fd_sc_hd__sdlclkp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdlclkp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 0.955000 1.195000 1.445000 ;
        RECT 0.855000 1.445000 1.240000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.570000 0.255000 6.840000 0.825000 ;
        RECT 6.570000 1.495000 6.840000 2.465000 ;
        RECT 6.670000 0.825000 6.840000 1.055000 ;
        RECT 6.670000 1.055000 7.275000 1.315000 ;
        RECT 6.670000 1.315000 6.840000 1.495000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.340000 1.665000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.705000 0.955000 6.050000 1.265000 ;
        RECT 4.705000 1.265000 4.925000 1.325000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.195000 0.785000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.515000  0.785000 0.685000 2.125000 ;
      RECT 0.515000  2.125000 1.260000 2.465000 ;
      RECT 1.015000  0.255000 1.195000 0.615000 ;
      RECT 1.365000  0.255000 2.500000 0.535000 ;
      RECT 1.365000  0.705000 1.705000 1.205000 ;
      RECT 1.365000  1.205000 1.865000 1.325000 ;
      RECT 1.410000  1.325000 1.865000 1.955000 ;
      RECT 1.430000  2.125000 2.205000 2.465000 ;
      RECT 1.875000  0.705000 2.160000 1.035000 ;
      RECT 2.035000  1.205000 3.015000 1.375000 ;
      RECT 2.035000  1.375000 2.205000 2.125000 ;
      RECT 2.330000  0.535000 2.500000 0.995000 ;
      RECT 2.330000  0.995000 3.015000 1.205000 ;
      RECT 2.375000  1.575000 2.545000 1.635000 ;
      RECT 2.375000  1.635000 3.405000 1.905000 ;
      RECT 2.375000  2.075000 3.015000 2.635000 ;
      RECT 2.670000  0.085000 3.015000 0.825000 ;
      RECT 3.185000  0.255000 3.405000 1.635000 ;
      RECT 3.185000  1.905000 3.405000 1.915000 ;
      RECT 3.185000  1.915000 5.490000 2.085000 ;
      RECT 3.185000  2.085000 3.405000 2.465000 ;
      RECT 3.575000  0.255000 3.925000 0.765000 ;
      RECT 3.575000  0.765000 4.000000 0.935000 ;
      RECT 3.575000  0.935000 3.745000 1.575000 ;
      RECT 3.575000  1.575000 4.040000 1.745000 ;
      RECT 3.575000  2.255000 5.530000 2.635000 ;
      RECT 3.915000  1.105000 4.460000 1.275000 ;
      RECT 4.095000  0.085000 4.425000 0.445000 ;
      RECT 4.170000  0.615000 4.825000 0.785000 ;
      RECT 4.170000  0.785000 4.460000 1.105000 ;
      RECT 4.210000  1.275000 4.460000 1.495000 ;
      RECT 4.210000  1.495000 5.010000 1.745000 ;
      RECT 4.595000  0.255000 4.825000 0.615000 ;
      RECT 5.100000  0.255000 5.310000 0.615000 ;
      RECT 5.100000  0.615000 6.400000 0.785000 ;
      RECT 5.180000  1.435000 5.650000 1.605000 ;
      RECT 5.180000  1.605000 5.490000 1.915000 ;
      RECT 5.490000  0.085000 6.400000 0.445000 ;
      RECT 5.700000  1.775000 6.400000 2.085000 ;
      RECT 5.700000  2.085000 5.870000 2.465000 ;
      RECT 5.820000  1.435000 6.400000 1.775000 ;
      RECT 6.070000  2.255000 6.400000 2.635000 ;
      RECT 6.230000  0.785000 6.400000 0.995000 ;
      RECT 6.230000  0.995000 6.500000 1.325000 ;
      RECT 6.230000  1.325000 6.400000 1.435000 ;
      RECT 7.010000  0.085000 7.275000 0.885000 ;
      RECT 7.010000  1.485000 7.275000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.530000  1.445000 1.700000 1.615000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 1.990000  0.765000 2.160000 0.935000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 3.830000  0.765000 4.000000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.290000  1.445000 4.460000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 1.470000 1.415000 1.760000 1.460000 ;
      RECT 1.470000 1.460000 4.520000 1.600000 ;
      RECT 1.470000 1.600000 1.760000 1.645000 ;
      RECT 1.930000 0.735000 2.220000 0.780000 ;
      RECT 1.930000 0.780000 4.060000 0.920000 ;
      RECT 1.930000 0.920000 2.220000 0.965000 ;
      RECT 3.770000 0.735000 4.060000 0.780000 ;
      RECT 3.770000 0.920000 4.060000 0.965000 ;
      RECT 4.230000 1.415000 4.520000 1.460000 ;
      RECT 4.230000 1.600000 4.520000 1.645000 ;
  END
END sky130_fd_sc_hd__sdlclkp_2
MACRO sky130_fd_sc_hd__sdlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.850000 0.955000 1.190000 1.325000 ;
        RECT 0.880000 1.325000 1.190000 1.445000 ;
        RECT 0.880000 1.445000 1.235000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.530000 0.255000 6.815000 0.825000 ;
        RECT 6.530000 1.495000 6.815000 2.465000 ;
        RECT 6.645000 0.825000 6.815000 1.495000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.340000 1.665000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.710000 0.955000 6.010000 1.265000 ;
        RECT 4.710000 1.265000 4.930000 1.325000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.190000 0.785000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.510000  0.785000 0.680000 1.460000 ;
      RECT 0.510000  1.460000 0.710000 1.755000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.540000  1.755000 0.710000 2.125000 ;
      RECT 0.540000  2.125000 1.255000 2.465000 ;
      RECT 1.015000  0.255000 1.190000 0.615000 ;
      RECT 1.360000  0.255000 2.495000 0.535000 ;
      RECT 1.360000  0.705000 1.700000 1.205000 ;
      RECT 1.360000  1.205000 1.860000 1.325000 ;
      RECT 1.405000  1.325000 1.860000 1.955000 ;
      RECT 1.425000  2.125000 2.200000 2.465000 ;
      RECT 1.870000  0.705000 2.155000 1.035000 ;
      RECT 2.030000  1.205000 3.010000 1.375000 ;
      RECT 2.030000  1.375000 2.200000 2.125000 ;
      RECT 2.325000  0.535000 2.495000 0.995000 ;
      RECT 2.325000  0.995000 3.010000 1.205000 ;
      RECT 2.370000  1.575000 2.540000 1.635000 ;
      RECT 2.370000  1.635000 3.400000 1.905000 ;
      RECT 2.370000  2.075000 3.010000 2.635000 ;
      RECT 2.665000  0.085000 3.010000 0.825000 ;
      RECT 3.180000  0.255000 3.400000 1.635000 ;
      RECT 3.180000  1.905000 3.400000 1.915000 ;
      RECT 3.180000  1.915000 5.450000 2.085000 ;
      RECT 3.180000  2.085000 3.400000 2.465000 ;
      RECT 3.580000  0.255000 3.910000 0.765000 ;
      RECT 3.580000  0.765000 4.005000 0.935000 ;
      RECT 3.580000  0.935000 3.750000 1.575000 ;
      RECT 3.580000  1.575000 3.990000 1.745000 ;
      RECT 3.580000  2.255000 5.490000 2.635000 ;
      RECT 3.920000  1.105000 4.465000 1.275000 ;
      RECT 4.080000  0.085000 4.410000 0.445000 ;
      RECT 4.160000  1.275000 4.465000 1.495000 ;
      RECT 4.160000  1.495000 4.960000 1.745000 ;
      RECT 4.175000  0.615000 4.830000 0.785000 ;
      RECT 4.175000  0.785000 4.465000 1.105000 ;
      RECT 4.580000  0.255000 4.830000 0.615000 ;
      RECT 5.010000  0.255000 5.270000 0.615000 ;
      RECT 5.010000  0.615000 6.360000 0.785000 ;
      RECT 5.140000  1.435000 5.610000 1.605000 ;
      RECT 5.140000  1.605000 5.450000 1.915000 ;
      RECT 5.505000  0.085000 6.360000 0.445000 ;
      RECT 5.660000  1.775000 6.360000 2.085000 ;
      RECT 5.660000  2.085000 5.830000 2.465000 ;
      RECT 5.780000  1.435000 6.360000 1.775000 ;
      RECT 6.030000  2.255000 6.360000 2.635000 ;
      RECT 6.190000  0.785000 6.360000 0.995000 ;
      RECT 6.190000  0.995000 6.460000 1.325000 ;
      RECT 6.190000  1.325000 6.360000 1.435000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  1.445000 1.695000 1.615000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  0.765000 2.155000 0.935000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 3.835000  0.765000 4.005000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.295000  1.445000 4.465000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.525000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 1.925000 0.735000 2.215000 0.780000 ;
      RECT 1.925000 0.780000 4.065000 0.920000 ;
      RECT 1.925000 0.920000 2.215000 0.965000 ;
      RECT 3.775000 0.735000 4.065000 0.780000 ;
      RECT 3.775000 0.920000 4.065000 0.965000 ;
      RECT 4.235000 1.415000 4.525000 1.460000 ;
      RECT 4.235000 1.600000 4.525000 1.645000 ;
  END
END sky130_fd_sc_hd__sdlclkp_1
MACRO sky130_fd_sc_hd__sdlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdlclkp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855000 0.955000 1.195000 1.445000 ;
        RECT 0.855000 1.445000 1.240000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.500000 0.255000 6.830000 0.445000 ;
        RECT 6.580000 0.445000 6.830000 0.715000 ;
        RECT 6.580000 0.715000 7.220000 0.885000 ;
        RECT 6.580000 1.485000 7.220000 1.655000 ;
        RECT 6.580000 1.655000 6.830000 2.465000 ;
        RECT 7.050000 0.885000 7.220000 1.055000 ;
        RECT 7.050000 1.055000 8.195000 1.315000 ;
        RECT 7.050000 1.315000 7.220000 1.485000 ;
        RECT 7.420000 0.255000 7.720000 1.055000 ;
        RECT 7.420000 1.315000 7.720000 2.465000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.345000 1.665000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.406500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.725000 0.995000 4.945000 1.325000 ;
      LAYER mcon ;
        RECT 4.770000 1.105000 4.940000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.685000 0.995000 6.065000 1.325000 ;
      LAYER mcon ;
        RECT 5.710000 1.105000 5.880000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.710000 1.075000 5.000000 1.120000 ;
        RECT 4.710000 1.120000 5.940000 1.260000 ;
        RECT 4.710000 1.260000 5.000000 1.305000 ;
        RECT 5.650000 1.075000 5.940000 1.120000 ;
        RECT 5.650000 1.260000 5.940000 1.305000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.195000 0.785000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.515000  0.785000 0.685000 2.125000 ;
      RECT 0.515000  2.125000 1.260000 2.465000 ;
      RECT 1.015000  0.255000 1.195000 0.615000 ;
      RECT 1.365000  0.255000 2.500000 0.535000 ;
      RECT 1.365000  0.705000 1.705000 1.205000 ;
      RECT 1.365000  1.205000 1.865000 1.325000 ;
      RECT 1.410000  1.325000 1.865000 1.955000 ;
      RECT 1.430000  2.125000 2.205000 2.465000 ;
      RECT 1.875000  0.705000 2.160000 1.035000 ;
      RECT 2.035000  1.205000 3.015000 1.375000 ;
      RECT 2.035000  1.375000 2.205000 2.125000 ;
      RECT 2.330000  0.535000 2.500000 0.995000 ;
      RECT 2.330000  0.995000 3.015000 1.205000 ;
      RECT 2.375000  1.575000 2.545000 1.635000 ;
      RECT 2.375000  1.635000 3.405000 1.905000 ;
      RECT 2.375000  2.075000 3.015000 2.635000 ;
      RECT 2.670000  0.085000 3.015000 0.825000 ;
      RECT 3.185000  0.255000 3.405000 1.635000 ;
      RECT 3.185000  1.905000 3.405000 1.915000 ;
      RECT 3.185000  1.915000 5.515000 2.085000 ;
      RECT 3.185000  2.085000 3.405000 2.465000 ;
      RECT 3.595000  0.255000 3.925000 0.765000 ;
      RECT 3.595000  0.765000 4.020000 0.935000 ;
      RECT 3.595000  0.935000 3.765000 1.575000 ;
      RECT 3.595000  1.575000 4.005000 1.745000 ;
      RECT 3.595000  2.255000 5.515000 2.635000 ;
      RECT 3.935000  1.105000 4.480000 1.275000 ;
      RECT 4.095000  0.085000 4.425000 0.445000 ;
      RECT 4.175000  1.275000 4.480000 1.495000 ;
      RECT 4.175000  1.495000 4.975000 1.745000 ;
      RECT 4.190000  0.615000 4.845000 0.785000 ;
      RECT 4.190000  0.785000 4.480000 1.105000 ;
      RECT 4.595000  0.255000 4.845000 0.615000 ;
      RECT 5.015000  0.255000 5.435000 0.615000 ;
      RECT 5.015000  0.615000 6.410000 0.785000 ;
      RECT 5.165000  0.995000 5.515000 1.915000 ;
      RECT 5.605000  0.085000 6.330000 0.445000 ;
      RECT 5.685000  1.495000 6.410000 2.085000 ;
      RECT 5.685000  2.085000 5.855000 2.465000 ;
      RECT 6.055000  2.255000 6.385000 2.635000 ;
      RECT 6.240000  0.785000 6.410000 1.055000 ;
      RECT 6.240000  1.055000 6.880000 1.315000 ;
      RECT 6.240000  1.315000 6.410000 1.495000 ;
      RECT 7.000000  0.085000 7.250000 0.545000 ;
      RECT 7.000000  1.825000 7.250000 2.635000 ;
      RECT 7.890000  0.085000 8.195000 0.885000 ;
      RECT 7.890000  1.485000 8.195000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.530000  1.445000 1.700000 1.615000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 1.990000  0.765000 2.160000 0.935000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 3.850000  0.765000 4.020000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.310000  1.445000 4.480000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 1.470000 1.415000 1.760000 1.460000 ;
      RECT 1.470000 1.460000 4.540000 1.600000 ;
      RECT 1.470000 1.600000 1.760000 1.645000 ;
      RECT 1.930000 0.735000 2.220000 0.780000 ;
      RECT 1.930000 0.780000 4.080000 0.920000 ;
      RECT 1.930000 0.920000 2.220000 0.965000 ;
      RECT 3.790000 0.735000 4.080000 0.780000 ;
      RECT 3.790000 0.920000 4.080000 0.965000 ;
      RECT 4.250000 1.415000 4.540000 1.460000 ;
      RECT 4.250000 1.600000 4.540000 1.645000 ;
  END
END sky130_fd_sc_hd__sdlclkp_4
MACRO sky130_fd_sc_hd__lpflow_inputiso1p_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso1p_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.765000 0.500000 1.325000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.765000 1.275000 1.325000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.509000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.255000 2.180000 0.825000 ;
        RECT 1.645000 1.845000 2.180000 2.465000 ;
        RECT 1.865000 0.825000 2.180000 1.845000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.250000  0.085000 0.490000 0.595000 ;
      RECT 0.270000  1.495000 1.695000 1.665000 ;
      RECT 0.270000  1.665000 0.660000 1.840000 ;
      RECT 0.670000  0.265000 0.950000 0.595000 ;
      RECT 0.670000  0.595000 0.840000 1.495000 ;
      RECT 1.145000  1.835000 1.475000 2.635000 ;
      RECT 1.180000  0.085000 1.395000 0.595000 ;
      RECT 1.525000  0.995000 1.695000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso1p_1
MACRO sky130_fd_sc_hd__tapvgnd2_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvgnd2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.315000 0.845000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.085000 1.755000 0.375000 1.985000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  1.470000 0.375000 2.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  1.785000 0.315000 1.955000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__tapvgnd2_1
MACRO sky130_fd_sc_hd__a22o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 0.675000 1.720000 1.075000 ;
        RECT 1.510000 1.075000 1.840000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.010000 1.075000 2.415000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765000 1.075000 1.240000 1.285000 ;
        RECT 1.020000 0.675000 1.240000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.575000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.900000 0.255000 3.160000 0.585000 ;
        RECT 2.900000 1.785000 3.160000 2.465000 ;
        RECT 2.990000 0.585000 3.160000 1.785000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  0.085000 0.545000 0.850000 ;
      RECT 0.095000  1.455000 2.815000 1.625000 ;
      RECT 0.095000  1.625000 0.425000 2.295000 ;
      RECT 0.095000  2.295000 1.265000 2.465000 ;
      RECT 0.595000  1.795000 2.230000 2.035000 ;
      RECT 0.595000  2.035000 0.825000 2.125000 ;
      RECT 0.820000  0.255000 2.145000 0.505000 ;
      RECT 0.935000  2.255000 1.265000 2.295000 ;
      RECT 1.455000  2.215000 1.810000 2.635000 ;
      RECT 1.975000  0.505000 2.145000 0.735000 ;
      RECT 1.975000  0.735000 2.815000 0.905000 ;
      RECT 1.980000  2.035000 2.230000 2.465000 ;
      RECT 2.355000  0.085000 2.685000 0.565000 ;
      RECT 2.400000  1.875000 2.730000 2.635000 ;
      RECT 2.645000  0.905000 2.815000 1.455000 ;
      RECT 3.330000  0.085000 3.500000 0.985000 ;
      RECT 3.330000  1.445000 3.500000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a22o_2
MACRO sky130_fd_sc_hd__a22o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.900000 1.075000 5.395000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.350000 1.075000 4.680000 1.445000 ;
        RECT 4.350000 1.445000 5.735000 1.615000 ;
        RECT 5.565000 1.075000 6.355000 1.275000 ;
        RECT 5.565000 1.275000 5.735000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.125000 1.075000 3.680000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.420000 1.075000 2.955000 1.445000 ;
        RECT 2.420000 1.445000 4.180000 1.615000 ;
        RECT 3.850000 1.075000 4.180000 1.445000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.725000 1.770000 0.905000 ;
        RECT 0.085000 0.905000 0.370000 1.445000 ;
        RECT 0.085000 1.445000 1.730000 1.615000 ;
        RECT 0.600000 0.265000 0.930000 0.725000 ;
        RECT 0.640000 1.615000 0.890000 2.465000 ;
        RECT 1.440000 0.255000 1.770000 0.725000 ;
        RECT 1.480000 1.615000 1.730000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.220000  1.825000 0.470000 2.635000 ;
      RECT 0.260000  0.085000 0.430000 0.555000 ;
      RECT 0.540000  1.075000 2.230000 1.275000 ;
      RECT 1.060000  1.795000 1.310000 2.635000 ;
      RECT 1.100000  0.085000 1.270000 0.555000 ;
      RECT 1.900000  1.275000 2.230000 1.785000 ;
      RECT 1.900000  1.785000 3.930000 1.955000 ;
      RECT 1.900000  2.125000 2.150000 2.635000 ;
      RECT 1.940000  0.085000 2.630000 0.555000 ;
      RECT 1.940000  0.735000 5.310000 0.905000 ;
      RECT 1.940000  0.905000 2.230000 1.075000 ;
      RECT 2.420000  2.125000 2.670000 2.295000 ;
      RECT 2.420000  2.295000 4.430000 2.465000 ;
      RECT 2.800000  0.255000 3.970000 0.475000 ;
      RECT 2.840000  1.955000 3.090000 2.125000 ;
      RECT 3.170000  0.645000 3.605000 0.735000 ;
      RECT 3.260000  2.125000 3.510000 2.295000 ;
      RECT 3.680000  1.955000 3.930000 2.125000 ;
      RECT 4.100000  1.785000 6.110000 1.955000 ;
      RECT 4.100000  1.955000 4.430000 2.295000 ;
      RECT 4.185000  0.085000 4.355000 0.555000 ;
      RECT 4.560000  0.255000 5.730000 0.475000 ;
      RECT 4.600000  2.125000 4.850000 2.635000 ;
      RECT 4.935000  0.645000 5.310000 0.735000 ;
      RECT 5.020000  1.955000 5.270000 2.465000 ;
      RECT 5.440000  2.125000 5.690000 2.635000 ;
      RECT 5.480000  0.475000 5.730000 0.895000 ;
      RECT 5.900000  0.085000 6.070000 0.895000 ;
      RECT 5.905000  1.455000 6.110000 1.785000 ;
      RECT 5.905000  1.955000 6.110000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__a22o_4
MACRO sky130_fd_sc_hd__a22o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 0.675000 1.695000 1.075000 ;
        RECT 1.485000 1.075000 1.815000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.040000 2.395000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765000 1.075000 1.240000 1.285000 ;
        RECT 1.020000 0.675000 1.240000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.575000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875000 0.255000 3.135000 0.585000 ;
        RECT 2.875000 1.785000 3.135000 2.465000 ;
        RECT 2.965000 0.585000 3.135000 1.785000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  0.085000 0.545000 0.850000 ;
      RECT 0.090000  1.455000 1.265000 1.515000 ;
      RECT 0.090000  1.515000 2.795000 1.625000 ;
      RECT 0.090000  1.625000 0.345000 2.245000 ;
      RECT 0.090000  2.245000 0.425000 2.465000 ;
      RECT 0.595000  1.795000 0.780000 1.885000 ;
      RECT 0.595000  1.885000 2.205000 2.085000 ;
      RECT 0.595000  2.085000 0.825000 2.125000 ;
      RECT 0.820000  0.255000 2.120000 0.465000 ;
      RECT 0.935000  1.625000 2.735000 1.685000 ;
      RECT 0.935000  1.685000 1.265000 1.715000 ;
      RECT 1.370000  1.875000 2.205000 1.885000 ;
      RECT 1.430000  2.255000 1.785000 2.635000 ;
      RECT 1.950000  0.465000 2.120000 0.615000 ;
      RECT 1.950000  0.615000 2.705000 0.740000 ;
      RECT 1.950000  0.740000 2.795000 0.785000 ;
      RECT 1.955000  2.085000 2.205000 2.465000 ;
      RECT 2.375000  0.085000 2.705000 0.445000 ;
      RECT 2.455000  1.855000 2.705000 2.635000 ;
      RECT 2.525000  0.785000 2.795000 0.905000 ;
      RECT 2.595000  1.480000 2.795000 1.515000 ;
      RECT 2.625000  0.905000 2.795000 1.480000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a22o_1
MACRO sky130_fd_sc_hd__clkinv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.576000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.065000 1.305000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.662600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.460000 1.755000 1.630000 ;
        RECT 0.155000 1.630000 0.410000 2.435000 ;
        RECT 1.010000 1.630000 1.270000 2.435000 ;
        RECT 1.025000 0.280000 1.250000 0.725000 ;
        RECT 1.025000 0.725000 1.755000 0.895000 ;
        RECT 1.475000 0.895000 1.755000 1.460000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.560000  0.085000 0.855000 0.610000 ;
      RECT 0.580000  1.800000 0.840000 2.635000 ;
      RECT 1.420000  0.085000 1.750000 0.555000 ;
      RECT 1.440000  1.800000 1.695000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinv_2
MACRO sky130_fd_sc_hd__clkinv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.152000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.065000 2.660000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.075200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.725000 3.135000 0.895000 ;
        RECT 0.105000 0.895000 0.275000 1.460000 ;
        RECT 0.105000 1.460000 3.135000 1.630000 ;
        RECT 0.605000 1.630000 0.860000 2.435000 ;
        RECT 1.030000 0.280000 1.290000 0.725000 ;
        RECT 1.465000 1.630000 1.720000 2.435000 ;
        RECT 1.890000 0.280000 2.145000 0.725000 ;
        RECT 2.320000 1.630000 2.580000 2.435000 ;
        RECT 2.835000 0.895000 3.135000 1.460000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.800000 0.430000 2.635000 ;
      RECT 0.565000  0.085000 0.860000 0.555000 ;
      RECT 1.030000  1.800000 1.290000 2.635000 ;
      RECT 1.460000  0.085000 1.720000 0.555000 ;
      RECT 1.890000  1.800000 2.150000 2.635000 ;
      RECT 2.315000  0.085000 2.615000 0.555000 ;
      RECT 2.750000  1.800000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinv_4
MACRO sky130_fd_sc_hd__clkinv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.375000 0.325000 1.325000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.336000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.840000 0.760000 ;
        RECT 0.515000 0.760000 1.295000 1.290000 ;
        RECT 0.515000 1.290000 0.845000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.085000  1.665000 0.345000 2.635000 ;
      RECT 1.010000  0.085000 1.295000 0.590000 ;
      RECT 1.015000  1.665000 1.295000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinv_1
MACRO sky130_fd_sc_hd__clkinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  4.608000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.345000 0.895000  2.155000 1.275000 ;
        RECT 8.930000 0.895000 10.710000 1.275000 ;
      LAYER mcon ;
        RECT 1.525000 1.105000 1.695000 1.275000 ;
        RECT 1.985000 1.105000 2.155000 1.275000 ;
        RECT 9.345000 1.105000 9.515000 1.275000 ;
        RECT 9.805000 1.105000 9.975000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465000 1.075000  2.215000 1.120000 ;
        RECT 1.465000 1.120000 10.035000 1.260000 ;
        RECT 1.465000 1.260000  2.215000 1.305000 ;
        RECT 9.285000 1.075000 10.035000 1.120000 ;
        RECT 9.285000 1.260000 10.035000 1.305000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.520900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.575000 1.455000 10.480000 1.665000 ;
        RECT  0.575000 1.665000  0.830000 2.465000 ;
        RECT  1.435000 1.665000  1.690000 2.450000 ;
        RECT  2.325000 0.280000  2.550000 1.415000 ;
        RECT  2.325000 1.415000  8.755000 1.455000 ;
        RECT  2.325000 1.665000  2.550000 2.465000 ;
        RECT  3.155000 0.280000  3.410000 1.415000 ;
        RECT  3.155000 1.665000  3.410000 2.450000 ;
        RECT  4.015000 0.280000  4.255000 1.415000 ;
        RECT  4.015000 1.665000  4.255000 2.450000 ;
        RECT  4.905000 0.280000  5.255000 1.415000 ;
        RECT  4.905000 1.665000  5.280000 2.450000 ;
        RECT  5.925000 0.280000  6.175000 1.415000 ;
        RECT  5.925000 1.665000  6.175000 2.450000 ;
        RECT  6.785000 0.280000  7.035000 1.415000 ;
        RECT  6.785000 1.665000  7.035000 2.450000 ;
        RECT  7.645000 0.280000  7.895000 1.415000 ;
        RECT  7.645000 1.665000  7.895000 2.450000 ;
        RECT  8.505000 0.280000  8.755000 1.415000 ;
        RECT  8.505000 1.665000  8.755000 2.450000 ;
        RECT  9.365000 1.665000  9.605000 2.450000 ;
        RECT 10.225000 1.665000 10.480000 2.450000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.140000  1.495000  0.405000 2.635000 ;
      RECT  1.000000  1.835000  1.260000 2.635000 ;
      RECT  1.855000  0.085000  2.125000 0.610000 ;
      RECT  1.865000  1.835000  2.120000 2.635000 ;
      RECT  2.720000  0.085000  2.985000 0.610000 ;
      RECT  2.720000  1.835000  2.980000 2.635000 ;
      RECT  3.580000  0.085000  3.845000 0.610000 ;
      RECT  3.585000  1.835000  3.840000 2.635000 ;
      RECT  4.465000  0.085000  4.730000 0.610000 ;
      RECT  4.465000  1.835000  4.720000 2.635000 ;
      RECT  5.490000  0.085000  5.755000 0.610000 ;
      RECT  5.490000  1.835000  5.745000 2.120000 ;
      RECT  5.490000  2.120000  5.750000 2.635000 ;
      RECT  6.350000  0.085000  6.575000 0.610000 ;
      RECT  6.355000  1.835000  6.610000 2.635000 ;
      RECT  7.210000  0.085000  7.475000 0.610000 ;
      RECT  7.215000  1.835000  7.470000 2.635000 ;
      RECT  8.070000  0.085000  8.335000 0.610000 ;
      RECT  8.075000  1.835000  8.330000 2.635000 ;
      RECT  8.930000  0.085000  9.195000 0.610000 ;
      RECT  8.935000  1.835000  9.190000 2.635000 ;
      RECT  9.795000  1.835000 10.050000 2.635000 ;
      RECT 10.650000  1.835000 10.910000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinv_16
MACRO sky130_fd_sc_hd__clkinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.304000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.035000 4.865000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.090400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.695000 5.440000 0.865000 ;
        RECT 0.115000 0.865000 0.285000 1.460000 ;
        RECT 0.115000 1.460000 5.440000 1.630000 ;
        RECT 0.565000 1.630000 0.805000 2.435000 ;
        RECT 1.405000 1.630000 1.645000 2.435000 ;
        RECT 1.535000 0.280000 1.725000 0.695000 ;
        RECT 2.245000 1.630000 2.495000 2.435000 ;
        RECT 2.395000 0.280000 2.585000 0.695000 ;
        RECT 3.080000 1.630000 3.325000 2.435000 ;
        RECT 3.255000 0.280000 3.445000 0.695000 ;
        RECT 3.920000 1.630000 4.175000 2.435000 ;
        RECT 4.115000 0.280000 4.305000 0.695000 ;
        RECT 4.765000 1.630000 5.005000 2.435000 ;
        RECT 5.170000 0.865000 5.440000 1.460000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.135000  1.800000 0.395000 2.635000 ;
      RECT 0.975000  1.800000 1.235000 2.635000 ;
      RECT 1.035000  0.085000 1.365000 0.525000 ;
      RECT 1.815000  1.800000 2.075000 2.635000 ;
      RECT 1.895000  0.085000 2.225000 0.525000 ;
      RECT 2.665000  1.800000 2.910000 2.635000 ;
      RECT 2.755000  0.085000 3.085000 0.525000 ;
      RECT 3.495000  1.800000 3.750000 2.635000 ;
      RECT 3.615000  0.085000 3.945000 0.525000 ;
      RECT 4.345000  1.800000 4.595000 2.635000 ;
      RECT 4.475000  0.085000 4.805000 0.525000 ;
      RECT 5.175000  1.800000 5.430000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__clkinv_8
MACRO sky130_fd_sc_hd__a311o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.945000 1.075000 7.275000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.255000 1.075000 6.040000 1.285000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.515000 1.075000 4.945000 1.285000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.075000 1.505000 1.285000 ;
        RECT 1.060000 1.285000 1.255000 1.625000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.745000 0.350000 1.625000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.904000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195000 0.295000 2.545000 0.465000 ;
        RECT 2.295000 0.465000 2.465000 0.715000 ;
        RECT 2.295000 0.715000 3.305000 0.885000 ;
        RECT 2.715000 1.545000 3.885000 1.715000 ;
        RECT 2.910000 0.885000 3.105000 1.545000 ;
        RECT 3.055000 0.295000 3.385000 0.465000 ;
        RECT 3.135000 0.465000 3.305000 0.715000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.095000  0.085000 0.345000 0.565000 ;
      RECT 0.175000  1.795000 0.345000 2.295000 ;
      RECT 0.175000  2.295000 2.025000 2.465000 ;
      RECT 0.515000  0.295000 0.845000 0.465000 ;
      RECT 0.515000  1.955000 0.845000 2.125000 ;
      RECT 0.595000  0.465000 0.765000 0.715000 ;
      RECT 0.595000  0.715000 2.025000 0.885000 ;
      RECT 0.595000  0.885000 0.765000 1.955000 ;
      RECT 1.015000  0.085000 1.185000 0.545000 ;
      RECT 1.015000  1.795000 1.185000 2.295000 ;
      RECT 1.355000  0.295000 1.685000 0.465000 ;
      RECT 1.435000  0.465000 1.605000 0.715000 ;
      RECT 1.435000  1.455000 2.385000 1.625000 ;
      RECT 1.435000  1.625000 1.605000 2.125000 ;
      RECT 1.855000  0.085000 2.025000 0.545000 ;
      RECT 1.855000  0.885000 2.025000 1.075000 ;
      RECT 1.855000  1.075000 2.705000 1.245000 ;
      RECT 1.855000  1.795000 2.025000 2.295000 ;
      RECT 2.195000  1.625000 2.385000 1.915000 ;
      RECT 2.195000  1.915000 6.765000 2.085000 ;
      RECT 2.295000  2.255000 2.625000 2.635000 ;
      RECT 2.715000  0.085000 2.885000 0.545000 ;
      RECT 3.135000  2.255000 3.465000 2.635000 ;
      RECT 3.275000  1.075000 4.320000 1.245000 ;
      RECT 3.555000  0.085000 4.065000 0.545000 ;
      RECT 3.975000  2.255000 4.305000 2.635000 ;
      RECT 4.150000  1.245000 4.320000 1.455000 ;
      RECT 4.150000  1.455000 6.685000 1.625000 ;
      RECT 4.275000  0.295000 4.605000 0.465000 ;
      RECT 4.355000  0.465000 4.525000 0.715000 ;
      RECT 4.355000  0.715000 6.005000 0.885000 ;
      RECT 4.475000  1.795000 4.645000 1.915000 ;
      RECT 4.475000  2.085000 4.645000 2.465000 ;
      RECT 4.775000  0.085000 4.945000 0.545000 ;
      RECT 4.815000  2.255000 5.175000 2.635000 ;
      RECT 5.255000  0.255000 7.270000 0.425000 ;
      RECT 5.255000  0.425000 6.345000 0.465000 ;
      RECT 5.375000  1.795000 5.545000 1.915000 ;
      RECT 5.375000  2.085000 5.545000 2.465000 ;
      RECT 5.675000  0.645000 6.005000 0.715000 ;
      RECT 5.715000  2.255000 6.045000 2.635000 ;
      RECT 6.175000  0.465000 6.345000 0.885000 ;
      RECT 6.515000  0.645000 6.845000 0.825000 ;
      RECT 6.515000  0.825000 6.685000 1.455000 ;
      RECT 6.595000  1.795000 6.765000 1.915000 ;
      RECT 6.595000  2.085000 6.765000 2.465000 ;
      RECT 6.935000  0.425000 7.270000 0.500000 ;
      RECT 6.935000  1.795000 7.270000 2.635000 ;
      RECT 7.015000  0.500000 7.270000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__a311o_4
MACRO sky130_fd_sc_hd__a311o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 0.765000 2.155000 0.995000 ;
        RECT 1.965000 0.995000 2.310000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 0.750000 1.705000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.905000 0.995000 1.240000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.620000 0.995000 3.095000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 0.995000 3.535000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.454000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.395000 0.670000 ;
        RECT 0.085000 0.670000 0.255000 1.785000 ;
        RECT 0.085000 1.785000 0.425000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.425000  0.995000 0.735000 1.325000 ;
      RECT 0.565000  0.655000 1.260000 0.825000 ;
      RECT 0.565000  0.825000 0.735000 0.995000 ;
      RECT 0.565000  1.325000 0.735000 1.495000 ;
      RECT 0.565000  1.495000 3.505000 1.665000 ;
      RECT 0.590000  0.085000 0.920000 0.465000 ;
      RECT 0.595000  2.175000 0.840000 2.635000 ;
      RECT 1.015000  1.835000 2.575000 2.005000 ;
      RECT 1.015000  2.005000 1.265000 2.465000 ;
      RECT 1.090000  0.255000 2.495000 0.425000 ;
      RECT 1.090000  0.425000 1.260000 0.655000 ;
      RECT 1.455000  2.255000 2.125000 2.635000 ;
      RECT 2.325000  0.425000 2.495000 0.655000 ;
      RECT 2.325000  0.655000 3.505000 0.825000 ;
      RECT 2.325000  2.005000 2.575000 2.465000 ;
      RECT 2.765000  0.085000 3.095000 0.485000 ;
      RECT 3.335000  0.255000 3.505000 0.655000 ;
      RECT 3.335000  1.665000 3.505000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a311o_1
MACRO sky130_fd_sc_hd__a311o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 0.605000 2.620000 0.995000 ;
        RECT 2.440000 0.995000 2.675000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 0.605000 2.165000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 0.995000 1.710000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895000 0.995000 3.235000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.695000 0.995000 4.005000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.295000 0.845000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.885000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 1.015000  0.085000 1.345000 0.465000 ;
      RECT 1.015000  0.655000 1.695000 0.825000 ;
      RECT 1.015000  0.825000 1.185000 1.495000 ;
      RECT 1.015000  1.495000 3.965000 1.665000 ;
      RECT 1.160000  1.835000 1.380000 2.635000 ;
      RECT 1.525000  0.255000 2.960000 0.425000 ;
      RECT 1.525000  0.425000 1.695000 0.655000 ;
      RECT 1.590000  1.835000 3.025000 2.005000 ;
      RECT 1.590000  2.005000 1.840000 2.465000 ;
      RECT 2.125000  2.255000 2.455000 2.635000 ;
      RECT 2.715000  2.005000 3.025000 2.465000 ;
      RECT 2.790000  0.425000 2.960000 0.655000 ;
      RECT 2.790000  0.655000 3.965000 0.825000 ;
      RECT 3.220000  0.085000 3.550000 0.485000 ;
      RECT 3.795000  0.255000 3.965000 0.655000 ;
      RECT 3.795000  1.665000 3.965000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a311o_2
MACRO sky130_fd_sc_hd__a32o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 0.665000 2.280000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.665000 1.800000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 0.995000 1.320000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.450000 0.660000 2.870000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.180000 0.995000 3.530000 1.325000 ;
        RECT 3.325000 1.325000 3.530000 1.615000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.544500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.300000 0.425000 0.560000 ;
        RECT 0.090000 0.560000 0.345000 1.915000 ;
        RECT 0.090000 1.915000 0.425000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.570000  0.995000 0.875000 1.325000 ;
      RECT 0.595000  0.085000 0.925000 0.485000 ;
      RECT 0.675000  1.835000 1.005000 2.635000 ;
      RECT 0.705000  0.655000 1.265000 0.825000 ;
      RECT 0.705000  0.825000 0.875000 0.995000 ;
      RECT 0.705000  1.325000 0.875000 1.495000 ;
      RECT 0.705000  1.495000 3.075000 1.665000 ;
      RECT 1.095000  0.315000 2.710000 0.485000 ;
      RECT 1.095000  0.485000 1.265000 0.655000 ;
      RECT 1.250000  1.875000 2.675000 2.045000 ;
      RECT 1.250000  2.045000 1.535000 2.465000 ;
      RECT 1.790000  2.215000 2.120000 2.635000 ;
      RECT 2.345000  2.045000 2.675000 2.295000 ;
      RECT 2.345000  2.295000 3.505000 2.465000 ;
      RECT 2.905000  1.665000 3.075000 2.125000 ;
      RECT 3.255000  0.085000 3.585000 0.805000 ;
      RECT 3.335000  1.795000 3.505000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a32o_1
MACRO sky130_fd_sc_hd__a32o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685000 0.955000 2.985000 1.325000 ;
        RECT 2.755000 0.415000 3.105000 0.610000 ;
        RECT 2.755000 0.610000 2.985000 0.955000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.165000 0.995000 3.545000 1.325000 ;
        RECT 3.305000 0.425000 3.545000 0.995000 ;
        RECT 3.305000 1.325000 3.545000 1.625000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 0.995000 4.055000 1.630000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.085000 1.075000 2.515000 1.245000 ;
        RECT 2.345000 1.245000 2.515000 1.445000 ;
        RECT 2.345000 1.445000 2.550000 1.615000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 0.745000 1.530000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.695500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.655000 0.845000 0.825000 ;
        RECT 0.135000 0.825000 0.345000 1.785000 ;
        RECT 0.135000 1.785000 1.185000 1.955000 ;
        RECT 0.135000 1.955000 0.345000 2.465000 ;
        RECT 1.015000 1.955000 1.185000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.465000 ;
      RECT 0.515000  2.125000 0.845000 2.635000 ;
      RECT 0.535000  0.995000 0.705000 1.445000 ;
      RECT 0.535000  1.445000 2.125000 1.615000 ;
      RECT 0.935000  0.085000 1.640000 0.445000 ;
      RECT 1.535000  1.785000 1.705000 2.295000 ;
      RECT 1.535000  2.295000 2.545000 2.465000 ;
      RECT 1.700000  0.615000 2.585000 0.785000 ;
      RECT 1.700000  0.785000 1.890000 1.445000 ;
      RECT 1.875000  1.615000 2.125000 1.945000 ;
      RECT 1.875000  1.945000 2.205000 2.115000 ;
      RECT 2.255000  0.275000 2.585000 0.615000 ;
      RECT 2.375000  1.795000 3.545000 1.965000 ;
      RECT 2.375000  1.965000 2.545000 2.295000 ;
      RECT 2.715000  2.140000 3.045000 2.635000 ;
      RECT 3.375000  1.965000 3.545000 2.465000 ;
      RECT 3.715000  0.085000 4.050000 0.805000 ;
      RECT 3.715000  1.915000 4.050000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a32o_2
MACRO sky130_fd_sc_hd__a32o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.280000 1.075000 5.075000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.335000 1.075000 4.030000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.075000 3.105000 1.295000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.630000 1.075000 6.780000 1.625000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.030000 1.075000 7.710000 1.295000 ;
        RECT 7.030000 1.295000 7.225000 1.635000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.635000 1.605000 0.805000 ;
        RECT 0.120000 0.805000 0.340000 1.495000 ;
        RECT 0.120000 1.495000 1.605000 1.665000 ;
        RECT 0.595000 0.255000 0.765000 0.635000 ;
        RECT 0.595000 1.665000 0.765000 2.465000 ;
        RECT 1.435000 0.255000 1.605000 0.635000 ;
        RECT 1.435000 1.665000 1.605000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.095000  1.915000 0.425000 2.635000 ;
      RECT 0.570000  0.995000 1.970000 1.325000 ;
      RECT 0.935000  0.085000 1.265000 0.465000 ;
      RECT 0.935000  1.915000 1.265000 2.635000 ;
      RECT 1.775000  0.085000 2.105000 0.465000 ;
      RECT 1.775000  1.915000 2.105000 2.635000 ;
      RECT 1.800000  1.325000 1.970000 1.495000 ;
      RECT 1.800000  1.495000 5.450000 1.665000 ;
      RECT 2.275000  0.255000 2.445000 0.655000 ;
      RECT 2.275000  0.655000 3.885000 0.825000 ;
      RECT 2.275000  1.915000 5.065000 2.085000 ;
      RECT 2.275000  2.085000 2.445000 2.465000 ;
      RECT 2.615000  0.085000 2.945000 0.465000 ;
      RECT 2.615000  2.255000 2.945000 2.635000 ;
      RECT 3.135000  0.295000 5.145000 0.465000 ;
      RECT 3.215000  2.085000 3.385000 2.465000 ;
      RECT 3.555000  2.255000 3.885000 2.635000 ;
      RECT 4.055000  2.085000 4.225000 2.465000 ;
      RECT 4.395000  0.635000 6.425000 0.805000 ;
      RECT 4.395000  2.255000 4.725000 2.635000 ;
      RECT 4.895000  2.085000 5.065000 2.255000 ;
      RECT 4.895000  2.255000 7.725000 2.425000 ;
      RECT 5.280000  0.805000 5.450000 1.495000 ;
      RECT 5.280000  1.665000 5.450000 1.905000 ;
      RECT 5.280000  1.905000 6.200000 1.915000 ;
      RECT 5.280000  1.915000 7.305000 2.075000 ;
      RECT 5.670000  0.295000 6.805000 0.465000 ;
      RECT 6.135000  2.075000 7.305000 2.085000 ;
      RECT 6.635000  0.255000 6.805000 0.295000 ;
      RECT 6.635000  0.465000 6.805000 0.645000 ;
      RECT 6.635000  0.645000 7.645000 0.815000 ;
      RECT 6.975000  0.085000 7.305000 0.465000 ;
      RECT 7.475000  0.255000 7.645000 0.645000 ;
      RECT 7.475000  1.755000 7.725000 2.255000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__a32o_4
MACRO sky130_fd_sc_hd__o31ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.440000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.075000 1.055000 2.465000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 1.075000 1.700000 1.325000 ;
        RECT 1.460000 1.325000 1.700000 2.405000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.330000 0.995000 2.675000 1.325000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.006000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 0.260000 2.675000 0.825000 ;
        RECT 1.945000 0.825000 2.160000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  1.495000 0.440000 2.635000 ;
      RECT 0.175000  0.085000 0.345000 0.905000 ;
      RECT 0.515000  0.255000 0.845000 0.735000 ;
      RECT 0.515000  0.735000 1.700000 0.905000 ;
      RECT 1.015000  0.085000 1.185000 0.565000 ;
      RECT 1.370000  0.255000 1.700000 0.735000 ;
      RECT 2.330000  1.495000 2.675000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__o31ai_1
MACRO sky130_fd_sc_hd__o31ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.055000 1.240000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.410000 1.055000 2.220000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.390000 1.055000 3.205000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 0.755000 4.515000 1.325000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.063500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335000 1.495000 4.515000 1.665000 ;
        RECT 2.335000 1.665000 2.665000 2.125000 ;
        RECT 3.175000 1.665000 3.505000 2.465000 ;
        RECT 3.675000 0.595000 4.005000 1.495000 ;
        RECT 4.175000 1.665000 4.515000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.255000 0.445000 0.715000 ;
      RECT 0.090000  0.715000 3.505000 0.885000 ;
      RECT 0.090000  1.495000 2.125000 1.665000 ;
      RECT 0.090000  1.665000 0.445000 2.465000 ;
      RECT 0.615000  0.085000 0.785000 0.545000 ;
      RECT 0.615000  1.835000 0.785000 2.635000 ;
      RECT 0.955000  0.255000 1.285000 0.715000 ;
      RECT 0.955000  1.665000 1.285000 2.465000 ;
      RECT 1.455000  0.085000 1.965000 0.545000 ;
      RECT 1.455000  1.835000 1.625000 2.295000 ;
      RECT 1.455000  2.295000 3.005000 2.465000 ;
      RECT 1.795000  1.665000 2.125000 2.125000 ;
      RECT 2.175000  0.255000 2.505000 0.715000 ;
      RECT 2.675000  0.085000 3.005000 0.545000 ;
      RECT 2.835000  1.835000 3.005000 2.295000 ;
      RECT 3.175000  0.255000 4.515000 0.425000 ;
      RECT 3.175000  0.425000 3.505000 0.715000 ;
      RECT 3.675000  1.835000 4.005000 2.635000 ;
      RECT 4.175000  0.425000 4.515000 0.585000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__o31ai_2
MACRO sky130_fd_sc_hd__o31ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.055000 1.780000 1.425000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.950000 1.055000 3.605000 1.425000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775000 1.055000 5.940000 1.275000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465000 1.055000 7.735000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.683800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775000 1.445000 7.735000 1.695000 ;
        RECT 5.770000 1.695000 5.940000 2.465000 ;
        RECT 6.110000 0.645000 7.280000 0.885000 ;
        RECT 6.110000 0.885000 6.295000 1.445000 ;
        RECT 6.610000 1.695000 6.780000 2.465000 ;
        RECT 7.450000 1.695000 7.735000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.090000  0.255000 0.445000 0.715000 ;
      RECT 0.090000  0.715000 5.940000 0.885000 ;
      RECT 0.090000  1.595000 2.125000 1.895000 ;
      RECT 0.090000  1.895000 0.445000 2.465000 ;
      RECT 0.615000  0.085000 0.785000 0.545000 ;
      RECT 0.615000  2.065000 0.785000 2.635000 ;
      RECT 0.955000  0.255000 1.285000 0.715000 ;
      RECT 0.955000  1.895000 1.285000 2.465000 ;
      RECT 1.455000  0.085000 1.625000 0.545000 ;
      RECT 1.455000  2.065000 1.625000 2.635000 ;
      RECT 1.795000  0.255000 2.125000 0.715000 ;
      RECT 1.795000  1.895000 2.125000 2.205000 ;
      RECT 1.795000  2.205000 3.885000 2.465000 ;
      RECT 2.295000  0.085000 2.465000 0.545000 ;
      RECT 2.295000  1.595000 3.605000 1.765000 ;
      RECT 2.295000  1.765000 2.465000 2.035000 ;
      RECT 2.635000  0.255000 2.965000 0.715000 ;
      RECT 2.635000  1.935000 2.965000 2.205000 ;
      RECT 3.135000  0.085000 3.305000 0.545000 ;
      RECT 3.135000  1.765000 3.605000 1.865000 ;
      RECT 3.135000  1.865000 5.600000 2.035000 ;
      RECT 3.475000  0.255000 3.805000 0.715000 ;
      RECT 3.995000  0.085000 4.640000 0.545000 ;
      RECT 4.080000  2.035000 5.600000 2.465000 ;
      RECT 4.810000  0.395000 4.980000 0.715000 ;
      RECT 5.150000  0.085000 5.600000 0.545000 ;
      RECT 5.770000  0.255000 7.735000 0.475000 ;
      RECT 5.770000  0.475000 5.940000 0.715000 ;
      RECT 6.110000  1.890000 6.440000 2.635000 ;
      RECT 6.950000  1.890000 7.280000 2.635000 ;
      RECT 7.450000  0.475000 7.735000 0.885000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__o31ai_4
MACRO sky130_fd_sc_hd__a41oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.785000 1.075000 2.455000 1.295000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.665000 1.075000 3.365000 1.285000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.545000 1.075000 4.575000 1.295000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.755000 1.075000 5.895000 1.295000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.075000 1.555000 1.280000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.645000 2.295000 0.815000 ;
        RECT 0.145000 0.815000 0.315000 1.455000 ;
        RECT 0.145000 1.455000 1.455000 1.625000 ;
        RECT 0.685000 0.255000 0.855000 0.645000 ;
        RECT 1.125000 1.625000 1.455000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.185000  0.085000 0.515000 0.465000 ;
      RECT 0.785000  1.795000 0.955000 2.295000 ;
      RECT 0.785000  2.295000 1.795000 2.465000 ;
      RECT 1.025000  0.085000 1.375000 0.465000 ;
      RECT 1.545000  0.295000 2.635000 0.465000 ;
      RECT 1.625000  1.535000 5.760000 1.705000 ;
      RECT 1.625000  1.705000 1.795000 2.295000 ;
      RECT 1.965000  1.915000 2.295000 2.635000 ;
      RECT 2.465000  0.465000 2.635000 0.645000 ;
      RECT 2.465000  0.645000 3.555000 0.815000 ;
      RECT 2.465000  1.705000 2.635000 2.465000 ;
      RECT 2.805000  0.295000 4.495000 0.465000 ;
      RECT 2.805000  1.915000 3.135000 2.635000 ;
      RECT 3.325000  1.705000 3.495000 2.465000 ;
      RECT 3.745000  0.645000 5.675000 0.815000 ;
      RECT 3.755000  1.915000 4.425000 2.635000 ;
      RECT 4.665000  1.705000 4.835000 2.465000 ;
      RECT 5.005000  0.085000 5.335000 0.465000 ;
      RECT 5.005000  1.915000 5.335000 2.635000 ;
      RECT 5.505000  0.255000 5.675000 0.645000 ;
      RECT 5.505000  1.705000 5.675000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__a41oi_2
MACRO sky130_fd_sc_hd__a41oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385000 0.995000 4.205000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.405000 1.075000 6.315000 1.285000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.560000 1.075000 7.955000 1.300000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285000 1.075000 9.975000 1.280000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.745000 1.305000 ;
        RECT 0.105000 1.305000 0.325000 1.965000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.575000 2.155000 1.685000 ;
        RECT 0.515000 1.685000 1.685000 1.745000 ;
        RECT 0.515000 1.745000 0.845000 2.085000 ;
        RECT 0.595000 0.255000 0.765000 0.635000 ;
        RECT 0.595000 0.635000 4.015000 0.805000 ;
        RECT 1.350000 1.495000 2.155000 1.575000 ;
        RECT 1.350000 1.745000 1.685000 2.085000 ;
        RECT 1.435000 0.255000 1.605000 0.635000 ;
        RECT 1.935000 0.805000 2.155000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.090000  0.085000  0.425000 0.465000 ;
      RECT 0.090000  2.255000  2.335000 2.425000 ;
      RECT 0.935000  0.085000  1.265000 0.465000 ;
      RECT 1.775000  0.085000  2.105000 0.465000 ;
      RECT 2.165000  1.905000  3.515000 2.075000 ;
      RECT 2.165000  2.075000  2.335000 2.255000 ;
      RECT 2.165000  2.425000  2.335000 2.465000 ;
      RECT 2.425000  0.295000  6.115000 0.465000 ;
      RECT 2.505000  2.255000  3.175000 2.635000 ;
      RECT 3.345000  1.575000  9.945000 1.745000 ;
      RECT 3.345000  1.745000  3.515000 1.905000 ;
      RECT 3.345000  2.075000  3.515000 2.465000 ;
      RECT 3.685000  1.915000  4.015000 2.635000 ;
      RECT 4.185000  1.745000  4.355000 2.425000 ;
      RECT 4.525000  0.635000  7.895000 0.805000 ;
      RECT 4.620000  1.915000  4.950000 2.635000 ;
      RECT 5.120000  1.745000  5.290000 2.465000 ;
      RECT 5.495000  1.915000  6.165000 2.635000 ;
      RECT 6.305000  0.295000  8.235000 0.465000 ;
      RECT 6.385000  1.745000  6.555000 2.465000 ;
      RECT 6.725000  1.915000  7.055000 2.635000 ;
      RECT 7.225000  1.745000  7.395000 2.465000 ;
      RECT 7.565000  1.915000  7.895000 2.635000 ;
      RECT 8.065000  0.255000  8.235000 0.295000 ;
      RECT 8.065000  0.465000  8.235000 0.635000 ;
      RECT 8.065000  0.635000  9.915000 0.805000 ;
      RECT 8.065000  1.745000  8.235000 2.465000 ;
      RECT 8.405000  0.085000  8.735000 0.465000 ;
      RECT 8.405000  1.915000  8.735000 2.635000 ;
      RECT 8.905000  0.255000  9.075000 0.635000 ;
      RECT 8.905000  1.745000  9.075000 2.465000 ;
      RECT 9.245000  0.085000  9.575000 0.465000 ;
      RECT 9.245000  1.915000  9.575000 2.635000 ;
      RECT 9.745000  0.255000  9.915000 0.635000 ;
      RECT 9.775000  1.745000  9.945000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__a41oi_4
MACRO sky130_fd_sc_hd__a41oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.780000 0.995000 3.085000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.890000 0.755000 2.210000 1.665000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.470000 0.755000 1.710000 1.665000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 0.965000 1.250000 1.665000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.965000 0.780000 1.665000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.669500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.285000 0.345000 0.615000 ;
        RECT 0.090000 0.615000 1.290000 0.785000 ;
        RECT 0.090000 0.785000 0.360000 1.845000 ;
        RECT 0.090000 1.845000 0.425000 2.425000 ;
        RECT 1.120000 0.295000 3.015000 0.465000 ;
        RECT 1.120000 0.465000 1.290000 0.615000 ;
        RECT 2.685000 0.465000 3.015000 0.805000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.595000  1.845000 3.015000 2.015000 ;
      RECT 0.595000  2.015000 0.845000 2.465000 ;
      RECT 0.620000  0.085000 0.950000 0.445000 ;
      RECT 1.120000  2.195000 1.450000 2.635000 ;
      RECT 1.760000  2.015000 1.930000 2.465000 ;
      RECT 2.215000  2.195000 2.545000 2.635000 ;
      RECT 2.765000  2.015000 3.015000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a41oi_1
MACRO sky130_fd_sc_hd__o32a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 0.995000 1.715000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.995000 2.160000 1.615000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415000 0.995000 2.635000 1.615000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.695000 1.075000 4.055000 1.245000 ;
        RECT 3.725000 1.245000 4.055000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.910000 0.995000 3.155000 1.615000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.845000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.885000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 1.015000  0.995000 1.325000 1.785000 ;
      RECT 1.015000  1.785000 3.525000 1.955000 ;
      RECT 1.015000  2.125000 1.525000 2.635000 ;
      RECT 1.095000  0.085000 1.425000 0.825000 ;
      RECT 1.695000  0.255000 2.025000 0.655000 ;
      RECT 1.695000  0.655000 3.025000 0.825000 ;
      RECT 2.195000  0.085000 2.525000 0.485000 ;
      RECT 2.695000  0.255000 4.055000 0.425000 ;
      RECT 2.695000  0.425000 3.025000 0.655000 ;
      RECT 2.695000  1.955000 3.025000 2.465000 ;
      RECT 3.195000  0.595000 3.525000 0.825000 ;
      RECT 3.325000  0.825000 3.525000 1.785000 ;
      RECT 3.695000  0.425000 4.055000 0.905000 ;
      RECT 3.695000  1.495000 4.055000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o32a_2
MACRO sky130_fd_sc_hd__o32a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 0.995000 1.175000 1.075000 ;
        RECT 1.005000 1.075000 1.255000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.995000 1.810000 1.325000 ;
        RECT 1.485000 1.325000 1.810000 2.125000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.980000 0.995000 2.255000 1.660000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.320000 0.995000 3.595000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 0.995000 2.795000 1.660000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.504000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.595000 0.825000 ;
        RECT 0.085000 0.825000 0.260000 1.495000 ;
        RECT 0.085000 1.495000 0.470000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.445000  0.995000 0.635000 1.075000 ;
      RECT 0.445000  1.075000 0.810000 1.325000 ;
      RECT 0.640000  1.325000 0.810000 1.495000 ;
      RECT 0.640000  1.495000 1.315000 1.665000 ;
      RECT 0.685000  1.835000 0.975000 2.635000 ;
      RECT 0.765000  0.085000 0.935000 0.645000 ;
      RECT 1.140000  0.255000 1.470000 0.655000 ;
      RECT 1.140000  0.655000 2.540000 0.825000 ;
      RECT 1.145000  1.665000 1.315000 2.295000 ;
      RECT 1.145000  2.295000 2.510000 2.465000 ;
      RECT 1.645000  0.085000 1.975000 0.485000 ;
      RECT 2.180000  1.835000 3.135000 2.085000 ;
      RECT 2.180000  2.085000 2.510000 2.295000 ;
      RECT 2.210000  0.255000 3.595000 0.465000 ;
      RECT 2.210000  0.465000 2.540000 0.655000 ;
      RECT 2.710000  0.635000 3.135000 0.825000 ;
      RECT 2.965000  0.825000 3.135000 1.835000 ;
      RECT 3.305000  0.465000 3.595000 0.735000 ;
      RECT 3.305000  1.495000 3.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o32a_1
MACRO sky130_fd_sc_hd__o32a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 1.075000 0.780000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.075000 1.700000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.010000 1.075000 2.625000 1.275000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.870000 1.075000 4.230000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.790000 1.075000 5.260000 1.275000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.305000 0.255000 6.635000 0.715000 ;
        RECT 6.305000 0.715000 8.135000 0.905000 ;
        RECT 6.305000 1.495000 8.135000 1.665000 ;
        RECT 6.305000 1.665000 6.635000 2.465000 ;
        RECT 7.145000 0.255000 7.475000 0.715000 ;
        RECT 7.145000 1.665000 7.475000 2.465000 ;
        RECT 7.645000 0.905000 8.135000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 2.965000 0.885000 ;
      RECT 0.085000  1.445000 1.265000 1.665000 ;
      RECT 0.085000  1.665000 0.425000 2.465000 ;
      RECT 0.515000  0.085000 2.545000 0.465000 ;
      RECT 0.595000  1.835000 0.765000 2.635000 ;
      RECT 0.935000  1.665000 1.265000 2.295000 ;
      RECT 0.935000  2.295000 2.105000 2.465000 ;
      RECT 1.435000  1.445000 2.625000 1.690000 ;
      RECT 1.435000  1.690000 1.605000 2.045000 ;
      RECT 1.775000  1.860000 2.105000 2.295000 ;
      RECT 2.295000  1.690000 2.625000 2.295000 ;
      RECT 2.295000  2.295000 3.465000 2.465000 ;
      RECT 2.715000  0.255000 5.695000 0.465000 ;
      RECT 2.715000  0.465000 2.965000 0.635000 ;
      RECT 2.795000  1.105000 3.645000 1.275000 ;
      RECT 2.795000  1.275000 2.965000 2.045000 ;
      RECT 3.135000  1.445000 3.465000 2.295000 ;
      RECT 3.455000  0.635000 5.775000 0.805000 ;
      RECT 3.455000  0.805000 3.645000 1.105000 ;
      RECT 3.655000  1.445000 3.985000 1.785000 ;
      RECT 3.655000  1.785000 4.825000 1.955000 ;
      RECT 3.655000  1.955000 3.985000 2.465000 ;
      RECT 4.155000  2.125000 4.325000 2.635000 ;
      RECT 4.400000  0.805000 4.620000 1.445000 ;
      RECT 4.400000  1.445000 5.195000 1.615000 ;
      RECT 4.495000  1.955000 4.825000 2.285000 ;
      RECT 4.495000  2.285000 5.695000 2.465000 ;
      RECT 5.025000  1.615000 5.195000 2.115000 ;
      RECT 5.365000  1.445000 5.695000 2.285000 ;
      RECT 5.520000  0.805000 5.775000 1.075000 ;
      RECT 5.520000  1.075000 7.475000 1.245000 ;
      RECT 5.520000  1.245000 6.135000 1.265000 ;
      RECT 5.965000  0.085000 6.135000 0.885000 ;
      RECT 5.965000  1.835000 6.135000 2.635000 ;
      RECT 6.805000  0.085000 6.975000 0.545000 ;
      RECT 6.805000  1.835000 6.975000 2.635000 ;
      RECT 7.645000  0.085000 7.900000 0.545000 ;
      RECT 7.645000  1.835000 7.900000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
END sky130_fd_sc_hd__o32a_4
MACRO sky130_fd_sc_hd__dfrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855000 0.265000 9.105000 0.795000 ;
        RECT 8.855000 1.445000 9.105000 2.325000 ;
        RECT 8.900000 0.795000 9.105000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.090000  0.345000 0.345000 0.635000 ;
      RECT 0.090000  0.635000 0.840000 0.805000 ;
      RECT 0.090000  1.795000 0.840000 1.965000 ;
      RECT 0.090000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 2.465000 ;
      RECT 1.545000  0.085000 1.875000 0.445000 ;
      RECT 1.850000  2.175000 2.100000 2.635000 ;
      RECT 2.045000  0.305000 2.540000 0.475000 ;
      RECT 2.045000  0.475000 2.215000 1.835000 ;
      RECT 2.045000  1.835000 2.440000 2.005000 ;
      RECT 2.270000  2.005000 2.440000 2.135000 ;
      RECT 2.270000  2.135000 2.520000 2.465000 ;
      RECT 2.385000  0.765000 2.735000 1.385000 ;
      RECT 2.610000  1.575000 3.075000 1.965000 ;
      RECT 2.735000  2.135000 3.415000 2.465000 ;
      RECT 2.745000  0.305000 3.600000 0.475000 ;
      RECT 2.905000  0.765000 3.260000 0.985000 ;
      RECT 2.905000  0.985000 3.075000 1.575000 ;
      RECT 3.245000  1.185000 4.935000 1.355000 ;
      RECT 3.245000  1.355000 3.415000 2.135000 ;
      RECT 3.430000  0.475000 3.600000 1.185000 ;
      RECT 3.585000  1.865000 4.660000 2.035000 ;
      RECT 3.585000  2.035000 3.755000 2.375000 ;
      RECT 3.775000  1.525000 5.275000 1.695000 ;
      RECT 3.990000  2.205000 4.320000 2.635000 ;
      RECT 4.475000  0.085000 4.805000 0.545000 ;
      RECT 4.490000  2.035000 4.660000 2.375000 ;
      RECT 4.765000  1.005000 4.935000 1.185000 ;
      RECT 4.955000  2.175000 5.325000 2.635000 ;
      RECT 5.015000  0.275000 5.365000 0.445000 ;
      RECT 5.015000  0.445000 5.275000 0.835000 ;
      RECT 5.105000  0.835000 5.275000 1.525000 ;
      RECT 5.105000  1.695000 5.275000 1.835000 ;
      RECT 5.105000  1.835000 5.665000 2.005000 ;
      RECT 5.465000  0.705000 5.675000 1.495000 ;
      RECT 5.465000  1.495000 6.140000 1.655000 ;
      RECT 5.465000  1.655000 6.430000 1.665000 ;
      RECT 5.495000  2.005000 5.665000 2.465000 ;
      RECT 5.585000  0.255000 6.535000 0.535000 ;
      RECT 5.845000  0.705000 6.195000 1.325000 ;
      RECT 5.900000  2.125000 6.770000 2.465000 ;
      RECT 5.970000  1.665000 6.430000 1.955000 ;
      RECT 6.365000  0.535000 6.535000 1.315000 ;
      RECT 6.365000  1.315000 6.770000 1.485000 ;
      RECT 6.600000  1.485000 6.770000 1.575000 ;
      RECT 6.600000  1.575000 7.820000 1.745000 ;
      RECT 6.600000  1.745000 6.770000 2.125000 ;
      RECT 6.705000  0.085000 6.895000 0.525000 ;
      RECT 6.705000  0.695000 7.235000 0.865000 ;
      RECT 6.705000  0.865000 6.925000 1.145000 ;
      RECT 6.940000  2.175000 7.190000 2.635000 ;
      RECT 7.065000  0.295000 8.135000 0.465000 ;
      RECT 7.065000  0.465000 7.235000 0.695000 ;
      RECT 7.360000  1.915000 8.160000 2.085000 ;
      RECT 7.360000  2.085000 7.530000 2.375000 ;
      RECT 7.710000  2.255000 8.040000 2.635000 ;
      RECT 7.815000  0.465000 8.135000 0.820000 ;
      RECT 7.815000  0.820000 8.140000 0.995000 ;
      RECT 7.815000  0.995000 8.730000 1.295000 ;
      RECT 7.990000  1.295000 8.730000 1.325000 ;
      RECT 7.990000  1.325000 8.160000 1.915000 ;
      RECT 8.380000  0.085000 8.685000 0.545000 ;
      RECT 8.380000  1.495000 8.685000 2.635000 ;
      RECT 9.275000  0.085000 9.525000 0.840000 ;
      RECT 9.275000  1.495000 9.525000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.105000 0.780000 1.275000 ;
      RECT 1.015000  1.785000 1.185000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.105000 2.615000 1.275000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  1.785000 3.075000 1.955000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.025000  1.105000 6.195000 1.275000 ;
      RECT 6.025000  1.785000 6.195000 1.955000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.075000 0.840000 1.120000 ;
      RECT 0.550000 1.120000 6.255000 1.260000 ;
      RECT 0.550000 1.260000 0.840000 1.305000 ;
      RECT 0.955000 1.755000 1.245000 1.800000 ;
      RECT 0.955000 1.800000 6.255000 1.940000 ;
      RECT 0.955000 1.940000 1.245000 1.985000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrtp_2
MACRO sky130_fd_sc_hd__dfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  8.675000 0.255000  9.005000 0.735000 ;
        RECT  8.675000 0.735000 10.440000 0.905000 ;
        RECT  8.715000 1.455000 10.440000 1.625000 ;
        RECT  8.715000 1.625000  9.005000 2.465000 ;
        RECT  9.515000 0.255000  9.845000 0.735000 ;
        RECT  9.555000 1.625000  9.805000 2.465000 ;
        RECT 10.030000 0.905000 10.440000 1.455000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.770000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.090000  0.345000  0.345000 0.635000 ;
      RECT  0.090000  0.635000  0.840000 0.805000 ;
      RECT  0.090000  1.795000  0.840000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.545000  0.085000  1.875000 0.445000 ;
      RECT  1.850000  2.175000  2.100000 2.635000 ;
      RECT  2.045000  0.305000  2.540000 0.475000 ;
      RECT  2.045000  0.475000  2.215000 1.835000 ;
      RECT  2.045000  1.835000  2.440000 2.005000 ;
      RECT  2.270000  2.005000  2.440000 2.135000 ;
      RECT  2.270000  2.135000  2.520000 2.465000 ;
      RECT  2.385000  0.765000  2.735000 1.385000 ;
      RECT  2.610000  1.575000  3.075000 1.965000 ;
      RECT  2.735000  2.135000  3.415000 2.465000 ;
      RECT  2.745000  0.305000  3.600000 0.475000 ;
      RECT  2.905000  0.765000  3.260000 0.985000 ;
      RECT  2.905000  0.985000  3.075000 1.575000 ;
      RECT  3.245000  1.185000  4.935000 1.355000 ;
      RECT  3.245000  1.355000  3.415000 2.135000 ;
      RECT  3.430000  0.475000  3.600000 1.185000 ;
      RECT  3.585000  1.865000  4.660000 2.035000 ;
      RECT  3.585000  2.035000  3.755000 2.375000 ;
      RECT  3.775000  1.525000  5.275000 1.695000 ;
      RECT  3.990000  2.205000  4.320000 2.635000 ;
      RECT  4.475000  0.085000  4.805000 0.545000 ;
      RECT  4.490000  2.035000  4.660000 2.375000 ;
      RECT  4.765000  1.005000  4.935000 1.185000 ;
      RECT  4.955000  2.175000  5.325000 2.635000 ;
      RECT  5.015000  0.275000  5.365000 0.445000 ;
      RECT  5.015000  0.445000  5.275000 0.835000 ;
      RECT  5.105000  0.835000  5.275000 1.525000 ;
      RECT  5.105000  1.695000  5.275000 1.835000 ;
      RECT  5.105000  1.835000  5.665000 2.005000 ;
      RECT  5.465000  0.705000  5.675000 1.495000 ;
      RECT  5.465000  1.495000  6.140000 1.655000 ;
      RECT  5.465000  1.655000  6.430000 1.665000 ;
      RECT  5.495000  2.005000  5.665000 2.465000 ;
      RECT  5.585000  0.255000  6.535000 0.535000 ;
      RECT  5.845000  0.705000  6.195000 1.325000 ;
      RECT  5.900000  2.125000  6.770000 2.465000 ;
      RECT  5.970000  1.665000  6.430000 1.955000 ;
      RECT  6.365000  0.535000  6.535000 1.315000 ;
      RECT  6.365000  1.315000  6.770000 1.485000 ;
      RECT  6.600000  1.485000  6.770000 1.575000 ;
      RECT  6.600000  1.575000  7.820000 1.745000 ;
      RECT  6.600000  1.745000  6.770000 2.125000 ;
      RECT  6.705000  0.085000  6.895000 0.525000 ;
      RECT  6.705000  0.695000  7.235000 0.865000 ;
      RECT  6.705000  0.865000  6.925000 1.145000 ;
      RECT  6.940000  2.175000  7.190000 2.635000 ;
      RECT  7.065000  0.295000  8.135000 0.465000 ;
      RECT  7.065000  0.465000  7.235000 0.695000 ;
      RECT  7.360000  1.915000  8.160000 2.085000 ;
      RECT  7.360000  2.085000  7.530000 2.375000 ;
      RECT  7.710000  2.255000  8.040000 2.635000 ;
      RECT  7.815000  0.465000  8.135000 0.820000 ;
      RECT  7.815000  0.820000  8.140000 1.075000 ;
      RECT  7.815000  1.075000  9.845000 1.285000 ;
      RECT  7.815000  1.285000  8.160000 1.295000 ;
      RECT  7.990000  1.295000  8.160000 1.915000 ;
      RECT  8.335000  0.085000  8.505000 0.895000 ;
      RECT  8.335000  1.575000  8.505000 2.635000 ;
      RECT  9.175000  0.085000  9.345000 0.555000 ;
      RECT  9.175000  1.795000  9.345000 2.635000 ;
      RECT 10.015000  0.085000 10.185000 0.555000 ;
      RECT 10.015000  1.795000 10.185000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.610000  1.105000  0.780000 1.275000 ;
      RECT  1.015000  1.785000  1.185000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.105000  2.615000 1.275000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  1.785000  3.075000 1.955000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.025000  1.105000  6.195000 1.275000 ;
      RECT  6.025000  1.785000  6.195000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.075000 0.840000 1.120000 ;
      RECT 0.550000 1.120000 6.255000 1.260000 ;
      RECT 0.550000 1.260000 0.840000 1.305000 ;
      RECT 0.955000 1.755000 1.245000 1.800000 ;
      RECT 0.955000 1.800000 6.255000 1.940000 ;
      RECT 0.955000 1.940000 1.245000 1.985000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrtp_4
MACRO sky130_fd_sc_hd__dfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855000 0.265000 9.110000 0.795000 ;
        RECT 8.855000 1.445000 9.110000 2.325000 ;
        RECT 8.900000 0.795000 9.110000 1.445000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.090000  0.345000 0.345000 0.635000 ;
      RECT 0.090000  0.635000 0.840000 0.805000 ;
      RECT 0.090000  1.795000 0.840000 1.965000 ;
      RECT 0.090000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 2.465000 ;
      RECT 1.545000  0.085000 1.875000 0.445000 ;
      RECT 1.850000  2.175000 2.100000 2.635000 ;
      RECT 2.045000  0.305000 2.540000 0.475000 ;
      RECT 2.045000  0.475000 2.215000 1.835000 ;
      RECT 2.045000  1.835000 2.440000 2.005000 ;
      RECT 2.270000  2.005000 2.440000 2.135000 ;
      RECT 2.270000  2.135000 2.520000 2.465000 ;
      RECT 2.385000  0.765000 2.735000 1.385000 ;
      RECT 2.610000  1.575000 3.075000 1.965000 ;
      RECT 2.735000  2.135000 3.415000 2.465000 ;
      RECT 2.745000  0.305000 3.600000 0.475000 ;
      RECT 2.905000  0.765000 3.260000 0.985000 ;
      RECT 2.905000  0.985000 3.075000 1.575000 ;
      RECT 3.245000  1.185000 4.935000 1.355000 ;
      RECT 3.245000  1.355000 3.415000 2.135000 ;
      RECT 3.430000  0.475000 3.600000 1.185000 ;
      RECT 3.585000  1.865000 4.660000 2.035000 ;
      RECT 3.585000  2.035000 3.755000 2.375000 ;
      RECT 3.775000  1.525000 5.275000 1.695000 ;
      RECT 3.990000  2.205000 4.320000 2.635000 ;
      RECT 4.475000  0.085000 4.805000 0.545000 ;
      RECT 4.490000  2.035000 4.660000 2.375000 ;
      RECT 4.765000  1.005000 4.935000 1.185000 ;
      RECT 4.955000  2.175000 5.325000 2.635000 ;
      RECT 5.015000  0.275000 5.365000 0.445000 ;
      RECT 5.015000  0.445000 5.275000 0.835000 ;
      RECT 5.105000  0.835000 5.275000 1.525000 ;
      RECT 5.105000  1.695000 5.275000 1.835000 ;
      RECT 5.105000  1.835000 5.665000 2.005000 ;
      RECT 5.465000  0.705000 5.675000 1.495000 ;
      RECT 5.465000  1.495000 6.140000 1.655000 ;
      RECT 5.465000  1.655000 6.430000 1.665000 ;
      RECT 5.495000  2.005000 5.665000 2.465000 ;
      RECT 5.585000  0.255000 6.535000 0.535000 ;
      RECT 5.845000  0.705000 6.195000 1.325000 ;
      RECT 5.900000  2.125000 6.770000 2.465000 ;
      RECT 5.970000  1.665000 6.430000 1.955000 ;
      RECT 6.365000  0.535000 6.535000 1.315000 ;
      RECT 6.365000  1.315000 6.770000 1.485000 ;
      RECT 6.600000  1.485000 6.770000 1.575000 ;
      RECT 6.600000  1.575000 7.820000 1.745000 ;
      RECT 6.600000  1.745000 6.770000 2.125000 ;
      RECT 6.705000  0.085000 6.895000 0.525000 ;
      RECT 6.705000  0.695000 7.235000 0.865000 ;
      RECT 6.705000  0.865000 6.925000 1.145000 ;
      RECT 6.940000  2.175000 7.190000 2.635000 ;
      RECT 7.065000  0.295000 8.135000 0.465000 ;
      RECT 7.065000  0.465000 7.235000 0.695000 ;
      RECT 7.360000  1.915000 8.160000 2.085000 ;
      RECT 7.360000  2.085000 7.530000 2.375000 ;
      RECT 7.710000  2.255000 8.040000 2.635000 ;
      RECT 7.815000  0.465000 8.135000 0.820000 ;
      RECT 7.815000  0.820000 8.140000 0.995000 ;
      RECT 7.815000  0.995000 8.730000 1.295000 ;
      RECT 7.990000  1.295000 8.730000 1.325000 ;
      RECT 7.990000  1.325000 8.160000 1.915000 ;
      RECT 8.380000  0.085000 8.685000 0.545000 ;
      RECT 8.380000  1.495000 8.685000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.105000 0.780000 1.275000 ;
      RECT 1.015000  1.785000 1.185000 1.955000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.105000 2.615000 1.275000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  1.785000 3.075000 1.955000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.025000  1.105000 6.195000 1.275000 ;
      RECT 6.025000  1.785000 6.195000 1.955000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.075000 0.840000 1.120000 ;
      RECT 0.550000 1.120000 6.255000 1.260000 ;
      RECT 0.550000 1.260000 0.840000 1.305000 ;
      RECT 0.955000 1.755000 1.245000 1.800000 ;
      RECT 0.955000 1.800000 6.255000 1.940000 ;
      RECT 0.955000 1.940000 1.245000 1.985000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrtp_1
MACRO sky130_fd_sc_hd__mux4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.540000 0.375000 6.850000 0.995000 ;
        RECT 6.540000 0.995000 6.950000 1.075000 ;
        RECT 6.640000 1.075000 6.950000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.750000 0.715000 5.120000 1.395000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.840000 0.765000 1.240000 1.095000 ;
        RECT 1.025000 0.395000 1.240000 0.765000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.245000 0.715000 2.620000 1.015000 ;
        RECT 2.415000 1.015000 2.620000 1.320000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.393000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.975000 0.330000 1.745000 ;
      LAYER mcon ;
        RECT 0.150000 1.445000 0.320000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.010000 1.445000 1.395000 1.615000 ;
        RECT 1.225000 1.285000 1.395000 1.445000 ;
      LAYER mcon ;
        RECT 1.070000 1.445000 1.240000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.130000 1.245000 6.470000 1.645000 ;
      LAYER mcon ;
        RECT 6.130000 1.445000 6.300000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085000 1.415000 0.380000 1.460000 ;
        RECT 0.085000 1.460000 6.360000 1.600000 ;
        RECT 0.085000 1.600000 0.380000 1.645000 ;
        RECT 1.010000 1.415000 1.300000 1.460000 ;
        RECT 1.010000 1.600000 1.300000 1.645000 ;
        RECT 6.070000 1.415000 6.360000 1.460000 ;
        RECT 6.070000 1.600000 6.360000 1.645000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.303000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 0.715000 3.080000 1.320000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.360000 1.835000 7.770000 2.455000 ;
        RECT 7.440000 0.265000 7.770000 0.725000 ;
        RECT 7.460000 1.495000 7.770000 1.835000 ;
        RECT 7.600000 0.725000 7.770000 1.065000 ;
        RECT 7.600000 1.065000 8.685000 1.305000 ;
        RECT 7.600000 1.305000 7.770000 1.495000 ;
        RECT 8.360000 0.265000 8.685000 1.065000 ;
        RECT 8.360000 1.305000 8.685000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.135000  0.345000 0.345000 0.635000 ;
      RECT 0.135000  0.635000 0.670000 0.805000 ;
      RECT 0.135000  1.915000 1.905000 1.955000 ;
      RECT 0.135000  1.955000 0.670000 2.085000 ;
      RECT 0.135000  2.085000 0.345000 2.375000 ;
      RECT 0.500000  0.805000 0.670000 1.785000 ;
      RECT 0.500000  1.785000 1.905000 1.915000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 1.410000  0.705000 1.735000 1.035000 ;
      RECT 1.415000  2.125000 2.245000 2.295000 ;
      RECT 1.475000  0.365000 2.075000 0.535000 ;
      RECT 1.565000  1.035000 1.735000 1.575000 ;
      RECT 1.565000  1.575000 1.905000 1.785000 ;
      RECT 1.905000  0.535000 2.075000 1.235000 ;
      RECT 1.905000  1.235000 2.245000 1.405000 ;
      RECT 2.075000  1.405000 2.245000 2.125000 ;
      RECT 2.455000  0.085000 2.785000 0.545000 ;
      RECT 2.600000  2.055000 2.830000 2.635000 ;
      RECT 2.975000  1.785000 3.320000 1.955000 ;
      RECT 2.990000  0.295000 3.420000 0.465000 ;
      RECT 3.150000  1.490000 3.420000 1.660000 ;
      RECT 3.150000  1.660000 3.320000 1.785000 ;
      RECT 3.250000  0.465000 3.420000 1.060000 ;
      RECT 3.250000  1.060000 3.485000 1.390000 ;
      RECT 3.250000  1.390000 3.420000 1.490000 ;
      RECT 3.310000  2.125000 3.825000 2.295000 ;
      RECT 3.575000  1.810000 3.825000 2.125000 ;
      RECT 3.590000  0.345000 3.825000 0.675000 ;
      RECT 3.655000  0.675000 3.825000 1.810000 ;
      RECT 3.995000  0.345000 4.185000 2.125000 ;
      RECT 3.995000  2.125000 4.520000 2.295000 ;
      RECT 4.400000  0.255000 4.605000 0.585000 ;
      RECT 4.400000  0.585000 4.570000 1.565000 ;
      RECT 4.400000  1.565000 5.500000 1.735000 ;
      RECT 4.400000  1.735000 4.590000 1.895000 ;
      RECT 4.760000  2.005000 5.105000 2.635000 ;
      RECT 4.800000  0.085000 5.130000 0.545000 ;
      RECT 5.330000  0.295000 6.225000 0.465000 ;
      RECT 5.330000  0.465000 5.500000 1.565000 ;
      RECT 5.330000  1.735000 5.500000 2.155000 ;
      RECT 5.330000  2.155000 6.280000 2.325000 ;
      RECT 5.670000  0.705000 6.290000 1.035000 ;
      RECT 5.670000  1.035000 5.960000 1.985000 ;
      RECT 6.530000  2.125000 6.850000 2.295000 ;
      RECT 6.680000  1.495000 7.290000 1.665000 ;
      RECT 6.680000  1.665000 6.850000 2.125000 ;
      RECT 7.020000  0.085000 7.270000 0.815000 ;
      RECT 7.020000  1.835000 7.190000 2.635000 ;
      RECT 7.120000  0.995000 7.430000 1.325000 ;
      RECT 7.120000  1.325000 7.290000 1.495000 ;
      RECT 7.940000  0.085000 8.190000 0.885000 ;
      RECT 7.940000  1.495000 8.190000 2.635000 ;
      RECT 8.855000  0.085000 9.105000 0.885000 ;
      RECT 8.855000  1.495000 9.105000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.530000  1.785000 1.700000 1.955000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 1.990000  2.125000 2.160000 2.295000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.370000  2.125000 3.540000 2.295000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.290000  2.125000 4.460000 2.295000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.670000  1.785000 5.840000 1.955000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.590000  2.125000 6.760000 2.295000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 1.470000 1.755000 1.760000 1.800000 ;
      RECT 1.470000 1.800000 5.900000 1.940000 ;
      RECT 1.470000 1.940000 1.760000 1.985000 ;
      RECT 1.930000 2.095000 2.220000 2.140000 ;
      RECT 1.930000 2.140000 3.600000 2.280000 ;
      RECT 1.930000 2.280000 2.220000 2.325000 ;
      RECT 3.310000 2.095000 3.600000 2.140000 ;
      RECT 3.310000 2.280000 3.600000 2.325000 ;
      RECT 4.230000 2.095000 4.520000 2.140000 ;
      RECT 4.230000 2.140000 6.820000 2.280000 ;
      RECT 4.230000 2.280000 4.520000 2.325000 ;
      RECT 5.610000 1.755000 5.900000 1.800000 ;
      RECT 5.610000 1.940000 5.900000 1.985000 ;
      RECT 6.530000 2.095000 6.820000 2.140000 ;
      RECT 6.530000 2.280000 6.820000 2.325000 ;
  END
END sky130_fd_sc_hd__mux4_4
MACRO sky130_fd_sc_hd__mux4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 0.995000 1.240000 1.615000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.995000 0.495000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.250000 1.055000 5.580000 1.675000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.800000 1.055000 5.045000 1.675000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.265000 0.995000 3.565000 1.995000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055000 0.995000 6.345000 1.675000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.315000 0.255000 9.575000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.175000  0.260000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 1.185000 0.805000 ;
      RECT 0.175000  1.795000 1.705000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 1.015000  0.255000 2.090000 0.425000 ;
      RECT 1.015000  0.425000 1.185000 0.635000 ;
      RECT 1.015000  2.135000 1.185000 2.295000 ;
      RECT 1.015000  2.295000 2.545000 2.465000 ;
      RECT 1.410000  0.595000 1.750000 0.765000 ;
      RECT 1.410000  0.765000 1.700000 0.935000 ;
      RECT 1.410000  0.935000 1.580000 1.455000 ;
      RECT 1.410000  1.455000 2.045000 1.625000 ;
      RECT 1.535000  1.965000 1.705000 2.125000 ;
      RECT 1.875000  1.625000 2.045000 1.955000 ;
      RECT 1.875000  1.955000 2.205000 2.125000 ;
      RECT 1.920000  0.425000 2.090000 0.760000 ;
      RECT 2.080000  1.105000 2.620000 1.285000 ;
      RECT 2.260000  0.430000 2.620000 1.105000 ;
      RECT 2.260000  1.285000 2.620000 1.395000 ;
      RECT 2.260000  1.395000 3.065000 1.625000 ;
      RECT 2.375000  1.795000 2.545000 2.295000 ;
      RECT 2.715000  1.625000 3.065000 2.465000 ;
      RECT 2.800000  0.085000 3.090000 0.805000 ;
      RECT 3.235000  2.255000 3.565000 2.635000 ;
      RECT 3.380000  0.255000 4.980000 0.425000 ;
      RECT 3.380000  0.425000 3.550000 0.795000 ;
      RECT 3.720000  0.595000 4.050000 0.845000 ;
      RECT 3.735000  0.845000 4.050000 0.920000 ;
      RECT 3.735000  0.920000 3.905000 1.445000 ;
      RECT 3.735000  1.445000 4.495000 1.615000 ;
      RECT 3.825000  1.785000 3.995000 2.295000 ;
      RECT 3.825000  2.295000 4.835000 2.465000 ;
      RECT 4.075000  1.095000 4.405000 1.105000 ;
      RECT 4.075000  1.105000 4.460000 1.265000 ;
      RECT 4.165000  1.615000 4.495000 2.125000 ;
      RECT 4.220000  0.595000 4.390000 0.715000 ;
      RECT 4.220000  0.715000 5.740000 0.885000 ;
      RECT 4.220000  0.885000 4.390000 0.925000 ;
      RECT 4.290000  1.265000 4.460000 1.275000 ;
      RECT 4.625000  0.425000 4.980000 0.465000 ;
      RECT 4.665000  1.915000 5.730000 2.085000 ;
      RECT 4.665000  2.085000 4.835000 2.295000 ;
      RECT 5.060000  2.255000 5.390000 2.635000 ;
      RECT 5.150000  0.085000 5.320000 0.545000 ;
      RECT 5.495000  0.295000 5.740000 0.715000 ;
      RECT 5.560000  2.085000 5.730000 2.465000 ;
      RECT 5.980000  2.255000 6.330000 2.635000 ;
      RECT 6.010000  0.085000 6.340000 0.465000 ;
      RECT 6.500000  2.135000 6.685000 2.465000 ;
      RECT 6.510000  0.325000 6.685000 0.655000 ;
      RECT 6.515000  0.655000 6.685000 1.105000 ;
      RECT 6.515000  1.105000 6.805000 1.275000 ;
      RECT 6.515000  1.275000 6.685000 2.135000 ;
      RECT 6.980000  0.765000 7.220000 0.935000 ;
      RECT 6.980000  0.935000 7.150000 2.135000 ;
      RECT 6.980000  2.135000 7.190000 2.465000 ;
      RECT 7.030000  0.255000 7.200000 0.415000 ;
      RECT 7.030000  0.415000 7.560000 0.585000 ;
      RECT 7.360000  2.255000 7.690000 2.295000 ;
      RECT 7.360000  2.295000 8.645000 2.465000 ;
      RECT 7.390000  0.585000 7.560000 1.755000 ;
      RECT 7.390000  1.755000 8.175000 1.985000 ;
      RECT 7.730000  0.255000 8.725000 0.425000 ;
      RECT 7.730000  0.425000 7.900000 0.585000 ;
      RECT 7.845000  1.985000 8.175000 2.125000 ;
      RECT 7.970000  0.765000 8.385000 0.925000 ;
      RECT 7.970000  0.925000 8.380000 0.935000 ;
      RECT 8.190000  1.105000 8.645000 1.275000 ;
      RECT 8.210000  0.595000 8.385000 0.765000 ;
      RECT 8.475000  1.665000 9.125000 1.835000 ;
      RECT 8.475000  1.835000 8.645000 2.295000 ;
      RECT 8.555000  0.425000 8.725000 0.715000 ;
      RECT 8.555000  0.715000 9.125000 0.885000 ;
      RECT 8.815000  2.255000 9.145000 2.635000 ;
      RECT 8.895000  0.085000 9.065000 0.545000 ;
      RECT 8.955000  0.885000 9.125000 1.665000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.530000  0.765000 1.700000 0.935000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.450000  1.105000 2.620000 1.275000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.290000  1.105000 4.460000 1.275000 ;
      RECT 4.325000  1.785000 4.495000 1.955000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.635000  1.105000 6.805000 1.275000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.050000  0.765000 7.220000 0.935000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.555000  1.785000 7.725000 1.955000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.475000  1.105000 8.645000 1.275000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 1.470000 0.735000 1.760000 0.780000 ;
      RECT 1.470000 0.780000 8.200000 0.920000 ;
      RECT 1.470000 0.920000 1.760000 0.965000 ;
      RECT 2.390000 1.075000 2.680000 1.120000 ;
      RECT 2.390000 1.120000 4.520000 1.260000 ;
      RECT 2.390000 1.260000 2.680000 1.305000 ;
      RECT 4.230000 1.075000 4.520000 1.120000 ;
      RECT 4.230000 1.260000 4.520000 1.305000 ;
      RECT 4.265000 1.755000 4.555000 1.800000 ;
      RECT 4.265000 1.800000 7.785000 1.940000 ;
      RECT 4.265000 1.940000 4.555000 1.985000 ;
      RECT 6.575000 1.075000 6.865000 1.120000 ;
      RECT 6.575000 1.120000 8.705000 1.260000 ;
      RECT 6.575000 1.260000 6.865000 1.305000 ;
      RECT 6.990000 0.735000 7.280000 0.780000 ;
      RECT 6.990000 0.920000 7.280000 0.965000 ;
      RECT 7.495000 1.755000 7.785000 1.800000 ;
      RECT 7.495000 1.940000 7.785000 1.985000 ;
      RECT 7.910000 0.735000 8.200000 0.780000 ;
      RECT 7.910000 0.920000 8.200000 0.965000 ;
      RECT 8.415000 1.075000 8.705000 1.120000 ;
      RECT 8.415000 1.260000 8.705000 1.305000 ;
  END
END sky130_fd_sc_hd__mux4_1
MACRO sky130_fd_sc_hd__mux4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 0.375000 6.845000 0.995000 ;
        RECT 6.535000 0.995000 6.945000 1.075000 ;
        RECT 6.635000 1.075000 6.945000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.745000 0.715000 5.115000 1.395000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 0.765000 1.235000 1.095000 ;
        RECT 1.020000 0.395000 1.235000 0.765000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.240000 0.715000 2.615000 1.015000 ;
        RECT 2.410000 1.015000 2.615000 1.320000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.393000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.975000 0.325000 1.745000 ;
      LAYER mcon ;
        RECT 0.145000 1.445000 0.315000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.005000 1.445000 1.390000 1.615000 ;
        RECT 1.220000 1.285000 1.390000 1.445000 ;
      LAYER mcon ;
        RECT 1.065000 1.445000 1.235000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.125000 1.245000 6.465000 1.645000 ;
      LAYER mcon ;
        RECT 6.125000 1.445000 6.295000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085000 1.415000 0.375000 1.460000 ;
        RECT 0.085000 1.460000 6.355000 1.600000 ;
        RECT 0.085000 1.600000 0.375000 1.645000 ;
        RECT 1.005000 1.415000 1.295000 1.460000 ;
        RECT 1.005000 1.600000 1.295000 1.645000 ;
        RECT 6.065000 1.415000 6.355000 1.460000 ;
        RECT 6.065000 1.600000 6.355000 1.645000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.303000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 0.715000 3.075000 1.320000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.355000 1.835000 7.765000 2.455000 ;
        RECT 7.435000 0.265000 7.765000 0.725000 ;
        RECT 7.455000 1.495000 7.765000 1.835000 ;
        RECT 7.595000 0.725000 7.765000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.170000  0.345000 0.345000 0.635000 ;
      RECT 0.170000  0.635000 0.665000 0.805000 ;
      RECT 0.175000  1.915000 1.900000 1.955000 ;
      RECT 0.175000  1.955000 0.665000 2.085000 ;
      RECT 0.175000  2.085000 0.345000 2.375000 ;
      RECT 0.495000  0.805000 0.665000 1.785000 ;
      RECT 0.495000  1.785000 1.900000 1.915000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 1.405000  0.705000 1.730000 1.035000 ;
      RECT 1.410000  2.125000 2.240000 2.295000 ;
      RECT 1.470000  0.365000 2.070000 0.535000 ;
      RECT 1.560000  1.035000 1.730000 1.575000 ;
      RECT 1.560000  1.575000 1.900000 1.785000 ;
      RECT 1.900000  0.535000 2.070000 1.235000 ;
      RECT 1.900000  1.235000 2.240000 1.405000 ;
      RECT 2.070000  1.405000 2.240000 2.125000 ;
      RECT 2.450000  0.085000 2.780000 0.545000 ;
      RECT 2.595000  2.055000 2.825000 2.635000 ;
      RECT 2.970000  1.785000 3.315000 1.955000 ;
      RECT 2.985000  0.295000 3.415000 0.465000 ;
      RECT 3.145000  1.490000 3.415000 1.660000 ;
      RECT 3.145000  1.660000 3.315000 1.785000 ;
      RECT 3.245000  0.465000 3.415000 1.060000 ;
      RECT 3.245000  1.060000 3.480000 1.390000 ;
      RECT 3.245000  1.390000 3.415000 1.490000 ;
      RECT 3.305000  2.125000 3.820000 2.295000 ;
      RECT 3.565000  1.810000 3.820000 2.125000 ;
      RECT 3.585000  0.345000 3.820000 0.675000 ;
      RECT 3.650000  0.675000 3.820000 1.810000 ;
      RECT 3.990000  0.345000 4.180000 2.125000 ;
      RECT 3.990000  2.125000 4.515000 2.295000 ;
      RECT 4.395000  0.255000 4.600000 0.585000 ;
      RECT 4.395000  0.585000 4.565000 1.565000 ;
      RECT 4.395000  1.565000 5.495000 1.735000 ;
      RECT 4.395000  1.735000 4.585000 1.895000 ;
      RECT 4.755000  2.005000 5.100000 2.635000 ;
      RECT 4.795000  0.085000 5.125000 0.545000 ;
      RECT 5.325000  0.295000 6.220000 0.465000 ;
      RECT 5.325000  0.465000 5.495000 1.565000 ;
      RECT 5.325000  1.735000 5.495000 2.155000 ;
      RECT 5.325000  2.155000 6.275000 2.325000 ;
      RECT 5.665000  0.705000 6.285000 1.035000 ;
      RECT 5.665000  1.035000 5.955000 1.985000 ;
      RECT 6.525000  2.125000 6.845000 2.295000 ;
      RECT 6.675000  1.495000 7.285000 1.665000 ;
      RECT 6.675000  1.665000 6.845000 2.125000 ;
      RECT 7.015000  0.085000 7.265000 0.815000 ;
      RECT 7.015000  1.835000 7.185000 2.635000 ;
      RECT 7.115000  0.995000 7.425000 1.325000 ;
      RECT 7.115000  1.325000 7.285000 1.495000 ;
      RECT 7.935000  0.085000 8.190000 0.885000 ;
      RECT 7.935000  1.495000 8.185000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  1.785000 1.695000 1.955000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.125000 2.155000 2.295000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.125000 3.535000 2.295000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.125000 4.455000 2.295000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  1.785000 5.835000 1.955000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.125000 6.755000 2.295000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.755000 1.755000 1.800000 ;
      RECT 1.465000 1.800000 5.895000 1.940000 ;
      RECT 1.465000 1.940000 1.755000 1.985000 ;
      RECT 1.925000 2.095000 2.215000 2.140000 ;
      RECT 1.925000 2.140000 3.595000 2.280000 ;
      RECT 1.925000 2.280000 2.215000 2.325000 ;
      RECT 3.305000 2.095000 3.595000 2.140000 ;
      RECT 3.305000 2.280000 3.595000 2.325000 ;
      RECT 4.225000 2.095000 4.515000 2.140000 ;
      RECT 4.225000 2.140000 6.815000 2.280000 ;
      RECT 4.225000 2.280000 4.515000 2.325000 ;
      RECT 5.605000 1.755000 5.895000 1.800000 ;
      RECT 5.605000 1.940000 5.895000 1.985000 ;
      RECT 6.525000 2.095000 6.815000 2.140000 ;
      RECT 6.525000 2.280000 6.815000 2.325000 ;
  END
END sky130_fd_sc_hd__mux4_2
MACRO sky130_fd_sc_hd__buf_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_12 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 1.075000 1.660000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.673000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275000 0.255000 2.445000 0.735000 ;
        RECT 2.275000 0.735000 6.645000 0.905000 ;
        RECT 2.275000 1.445000 6.645000 1.615000 ;
        RECT 2.275000 1.615000 2.445000 2.465000 ;
        RECT 3.115000 0.255000 3.285000 0.735000 ;
        RECT 3.115000 1.615000 3.285000 2.465000 ;
        RECT 3.955000 0.255000 4.125000 0.735000 ;
        RECT 3.955000 1.615000 4.125000 2.465000 ;
        RECT 4.710000 0.905000 6.645000 1.445000 ;
        RECT 4.795000 0.255000 4.965000 0.735000 ;
        RECT 4.795000 1.615000 4.965000 2.465000 ;
        RECT 5.635000 0.255000 5.805000 0.735000 ;
        RECT 5.635000 1.615000 5.805000 2.465000 ;
        RECT 6.475000 0.255000 6.645000 0.735000 ;
        RECT 6.475000 1.615000 6.645000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.570000 -0.085000 0.740000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.565000 ;
      RECT 0.175000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  1.445000 2.015000 1.615000 ;
      RECT 0.515000  1.615000 0.845000 2.465000 ;
      RECT 0.595000  0.255000 0.765000 0.735000 ;
      RECT 0.595000  0.735000 2.015000 0.905000 ;
      RECT 0.935000  0.085000 1.265000 0.565000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.355000  1.615000 1.685000 2.465000 ;
      RECT 1.435000  0.260000 1.605000 0.735000 ;
      RECT 1.775000  0.085000 2.105000 0.565000 ;
      RECT 1.840000  0.905000 2.015000 1.075000 ;
      RECT 1.840000  1.075000 4.465000 1.245000 ;
      RECT 1.840000  1.245000 2.015000 1.445000 ;
      RECT 1.855000  1.835000 2.025000 2.635000 ;
      RECT 2.615000  0.085000 2.945000 0.565000 ;
      RECT 2.615000  1.835000 2.945000 2.635000 ;
      RECT 3.455000  0.085000 3.785000 0.565000 ;
      RECT 3.455000  1.835000 3.785000 2.635000 ;
      RECT 4.295000  0.085000 4.625000 0.565000 ;
      RECT 4.295000  1.835000 4.625000 2.635000 ;
      RECT 5.135000  0.085000 5.465000 0.565000 ;
      RECT 5.135000  1.835000 5.465000 2.635000 ;
      RECT 5.975000  0.085000 6.305000 0.565000 ;
      RECT 5.975000  1.835000 6.305000 2.635000 ;
      RECT 6.815000  0.085000 7.145000 0.885000 ;
      RECT 6.815000  1.485000 7.145000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_12
MACRO sky130_fd_sc_hd__buf_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_6 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.280000 1.075000 1.185000 1.315000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.336500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.255000 1.865000 0.735000 ;
        RECT 1.695000 0.735000 3.545000 0.905000 ;
        RECT 1.695000 1.445000 3.545000 1.615000 ;
        RECT 1.695000 1.615000 1.865000 2.465000 ;
        RECT 2.210000 0.905000 3.545000 1.445000 ;
        RECT 2.535000 0.255000 2.705000 0.735000 ;
        RECT 2.535000 1.615000 2.705000 2.465000 ;
        RECT 3.375000 0.255000 3.545000 0.735000 ;
        RECT 3.375000 1.615000 3.545000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.435000  0.085000 0.605000 0.565000 ;
      RECT 0.435000  1.485000 0.605000 2.635000 ;
      RECT 0.775000  0.255000 1.105000 0.735000 ;
      RECT 0.775000  0.735000 1.525000 0.905000 ;
      RECT 0.775000  1.485000 1.525000 1.655000 ;
      RECT 0.775000  1.655000 1.105000 2.465000 ;
      RECT 1.275000  0.085000 1.445000 0.565000 ;
      RECT 1.275000  1.835000 1.515000 2.635000 ;
      RECT 1.355000  0.905000 1.525000 1.075000 ;
      RECT 1.355000  1.075000 1.825000 1.245000 ;
      RECT 1.355000  1.245000 1.525000 1.485000 ;
      RECT 2.035000  0.085000 2.365000 0.565000 ;
      RECT 2.035000  1.835000 2.365000 2.635000 ;
      RECT 2.875000  0.085000 3.205000 0.565000 ;
      RECT 2.875000  1.835000 3.205000 2.635000 ;
      RECT 3.715000  0.085000 4.045000 0.885000 ;
      RECT 3.715000  1.485000 4.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_6
MACRO sky130_fd_sc_hd__buf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.196500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.985000 0.445000 1.355000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.560000 1.295000 2.465000 ;
        RECT 1.035000 0.255000 1.295000 0.760000 ;
        RECT 1.115000 0.760000 1.295000 1.560000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.165000  1.535000 0.840000 1.705000 ;
      RECT 0.165000  1.705000 0.345000 2.465000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.525000  0.085000 0.855000 0.465000 ;
      RECT 0.525000  1.875000 0.855000 2.635000 ;
      RECT 0.670000  0.805000 0.840000 1.060000 ;
      RECT 0.670000  1.060000 0.945000 1.390000 ;
      RECT 0.670000  1.390000 0.840000 1.535000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_1
MACRO sky130_fd_sc_hd__buf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.240000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.855000 0.255000 2.025000 0.735000 ;
        RECT 1.855000 0.735000 4.545000 0.905000 ;
        RECT 1.855000 1.445000 4.545000 1.615000 ;
        RECT 1.855000 1.615000 2.025000 2.465000 ;
        RECT 2.695000 0.255000 2.865000 0.735000 ;
        RECT 2.695000 1.615000 2.865000 2.465000 ;
        RECT 3.535000 0.255000 3.705000 0.735000 ;
        RECT 3.535000 1.615000 3.705000 2.465000 ;
        RECT 4.290000 0.905000 4.545000 1.445000 ;
        RECT 4.375000 0.255000 4.545000 0.735000 ;
        RECT 4.375000 1.615000 4.545000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.095000  1.445000 1.595000 1.615000 ;
      RECT 0.095000  1.615000 0.425000 2.465000 ;
      RECT 0.175000  0.255000 0.345000 0.735000 ;
      RECT 0.175000  0.735000 1.595000 0.905000 ;
      RECT 0.515000  0.085000 0.845000 0.565000 ;
      RECT 0.595000  1.835000 0.765000 2.635000 ;
      RECT 0.935000  1.615000 1.265000 2.465000 ;
      RECT 1.015000  0.260000 1.185000 0.735000 ;
      RECT 1.355000  0.085000 1.685000 0.565000 ;
      RECT 1.420000  0.905000 1.595000 1.075000 ;
      RECT 1.420000  1.075000 4.045000 1.245000 ;
      RECT 1.420000  1.245000 1.595000 1.445000 ;
      RECT 1.435000  1.835000 1.605000 2.635000 ;
      RECT 2.195000  0.085000 2.525000 0.565000 ;
      RECT 2.195000  1.835000 2.525000 2.635000 ;
      RECT 3.035000  0.085000 3.365000 0.565000 ;
      RECT 3.035000  1.835000 3.365000 2.635000 ;
      RECT 3.875000  0.085000 4.205000 0.565000 ;
      RECT 3.875000  1.835000 4.205000 2.635000 ;
      RECT 4.715000  0.085000 5.045000 0.885000 ;
      RECT 4.715000  1.485000 5.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_8
MACRO sky130_fd_sc_hd__buf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.470000 1.315000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 0.255000 1.185000 0.735000 ;
        RECT 1.015000 0.735000 2.025000 0.905000 ;
        RECT 1.015000 1.445000 2.025000 1.615000 ;
        RECT 1.015000 1.615000 1.185000 2.465000 ;
        RECT 1.530000 0.905000 2.025000 1.445000 ;
        RECT 1.855000 0.255000 2.025000 0.735000 ;
        RECT 1.855000 1.615000 2.025000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  1.485000 0.810000 1.655000 ;
      RECT 0.095000  1.655000 0.425000 2.465000 ;
      RECT 0.175000  0.255000 0.345000 0.735000 ;
      RECT 0.175000  0.735000 0.810000 0.905000 ;
      RECT 0.525000  0.085000 0.765000 0.565000 ;
      RECT 0.595000  1.835000 0.835000 2.635000 ;
      RECT 0.640000  0.905000 0.810000 1.075000 ;
      RECT 0.640000  1.075000 1.140000 1.245000 ;
      RECT 0.640000  1.245000 0.810000 1.485000 ;
      RECT 1.355000  0.085000 1.685000 0.565000 ;
      RECT 1.355000  1.835000 1.685000 2.635000 ;
      RECT 2.195000  0.085000 2.525000 0.885000 ;
      RECT 2.195000  1.485000 2.525000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_4
MACRO sky130_fd_sc_hd__buf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.485000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 2.485000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 0.255000  3.285000 0.260000 ;
        RECT 3.035000 0.260000  3.365000 0.735000 ;
        RECT 3.035000 0.735000 10.035000 0.905000 ;
        RECT 3.035000 1.445000 10.035000 1.615000 ;
        RECT 3.035000 1.615000  3.365000 2.465000 ;
        RECT 3.875000 0.260000  4.205000 0.735000 ;
        RECT 3.875000 1.615000  4.205000 2.465000 ;
        RECT 3.955000 0.255000  4.125000 0.260000 ;
        RECT 4.715000 0.260000  5.045000 0.735000 ;
        RECT 4.715000 1.615000  5.045000 2.465000 ;
        RECT 4.795000 0.255000  4.965000 0.260000 ;
        RECT 5.555000 0.260000  5.885000 0.735000 ;
        RECT 5.555000 1.615000  5.885000 2.465000 ;
        RECT 6.395000 0.260000  6.725000 0.735000 ;
        RECT 6.395000 1.615000  6.725000 2.465000 ;
        RECT 7.235000 0.260000  7.565000 0.735000 ;
        RECT 7.235000 1.615000  7.565000 2.465000 ;
        RECT 8.075000 0.260000  8.405000 0.735000 ;
        RECT 8.075000 1.615000  8.405000 2.465000 ;
        RECT 8.915000 0.260000  9.245000 0.735000 ;
        RECT 8.915000 1.615000  9.245000 2.465000 ;
        RECT 9.655000 0.905000 10.035000 1.445000 ;
        RECT 9.760000 0.365000 10.035000 0.735000 ;
        RECT 9.760000 1.615000 10.035000 2.360000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.175000  0.085000  0.345000 0.905000 ;
      RECT 0.175000  1.445000  0.345000 2.635000 ;
      RECT 0.515000  0.260000  0.845000 0.735000 ;
      RECT 0.515000  0.735000  2.865000 0.905000 ;
      RECT 0.515000  1.445000  2.865000 1.615000 ;
      RECT 0.515000  1.615000  0.845000 2.465000 ;
      RECT 1.015000  0.085000  1.185000 0.565000 ;
      RECT 1.015000  1.835000  1.185000 2.635000 ;
      RECT 1.355000  0.260000  1.685000 0.735000 ;
      RECT 1.355000  1.615000  1.685000 2.465000 ;
      RECT 1.855000  0.085000  2.025000 0.565000 ;
      RECT 1.855000  1.835000  2.025000 2.635000 ;
      RECT 2.195000  0.260000  2.525000 0.735000 ;
      RECT 2.195000  1.615000  2.525000 2.465000 ;
      RECT 2.690000  0.905000  2.865000 1.075000 ;
      RECT 2.690000  1.075000  9.410000 1.275000 ;
      RECT 2.690000  1.275000  2.865000 1.445000 ;
      RECT 2.695000  0.085000  2.865000 0.565000 ;
      RECT 2.695000  1.835000  2.865000 2.635000 ;
      RECT 3.535000  0.085000  3.705000 0.565000 ;
      RECT 3.535000  1.835000  3.705000 2.635000 ;
      RECT 4.375000  0.085000  4.545000 0.565000 ;
      RECT 4.375000  1.835000  4.545000 2.635000 ;
      RECT 5.215000  0.085000  5.385000 0.565000 ;
      RECT 5.215000  1.835000  5.385000 2.635000 ;
      RECT 6.055000  0.085000  6.225000 0.565000 ;
      RECT 6.055000  1.835000  6.225000 2.635000 ;
      RECT 6.895000  0.085000  7.065000 0.565000 ;
      RECT 6.895000  1.835000  7.065000 2.635000 ;
      RECT 7.735000  0.085000  7.905000 0.565000 ;
      RECT 7.735000  1.835000  7.905000 2.635000 ;
      RECT 8.575000  0.085000  8.745000 0.565000 ;
      RECT 8.575000  1.835000  8.745000 2.635000 ;
      RECT 9.415000  0.085000  9.585000 0.565000 ;
      RECT 9.415000  1.835000  9.585000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_16
MACRO sky130_fd_sc_hd__buf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.440000 1.355000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.255000 1.315000 0.830000 ;
        RECT 1.060000 1.560000 1.315000 2.465000 ;
        RECT 1.145000 0.830000 1.315000 1.560000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.890000 0.805000 ;
      RECT 0.175000  1.535000 0.890000 1.705000 ;
      RECT 0.175000  1.705000 0.345000 2.465000 ;
      RECT 0.560000  0.085000 0.890000 0.465000 ;
      RECT 0.560000  1.875000 0.890000 2.635000 ;
      RECT 0.720000  0.805000 0.890000 0.995000 ;
      RECT 0.720000  0.995000 0.975000 1.325000 ;
      RECT 0.720000  1.325000 0.890000 1.535000 ;
      RECT 1.490000  0.085000 1.750000 0.925000 ;
      RECT 1.490000  1.485000 1.750000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_2
MACRO sky130_fd_sc_hd__xnor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.505000 1.075000 7.915000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.685000 0.995000 6.855000 1.445000 ;
        RECT 6.685000 1.445000 7.265000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.075000 2.640000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.350000 0.805000 0.925000 ;
        RECT 0.545000 0.925000 0.790000 1.440000 ;
        RECT 0.545000 1.440000 0.825000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.735000 ;
      RECT 0.085000  1.490000 0.375000 2.635000 ;
      RECT 0.960000  0.995000 1.165000 1.325000 ;
      RECT 0.975000  0.085000 1.225000 0.525000 ;
      RECT 0.990000  0.695000 1.565000 0.865000 ;
      RECT 0.990000  0.865000 1.165000 0.995000 ;
      RECT 0.995000  1.325000 1.165000 1.875000 ;
      RECT 0.995000  1.875000 1.680000 2.045000 ;
      RECT 0.995000  2.215000 1.330000 2.635000 ;
      RECT 1.395000  0.255000 2.965000 0.425000 ;
      RECT 1.395000  0.425000 1.565000 0.695000 ;
      RECT 1.395000  1.535000 2.980000 1.705000 ;
      RECT 1.510000  2.045000 1.680000 2.235000 ;
      RECT 1.510000  2.235000 2.980000 2.405000 ;
      RECT 1.735000  0.595000 1.905000 1.535000 ;
      RECT 2.020000  1.895000 4.520000 2.065000 ;
      RECT 2.205000  0.625000 3.425000 0.795000 ;
      RECT 2.205000  0.795000 2.585000 0.905000 ;
      RECT 2.530000  0.425000 2.965000 0.455000 ;
      RECT 2.810000  0.995000 3.085000 1.325000 ;
      RECT 2.810000  1.325000 2.980000 1.535000 ;
      RECT 3.135000  0.285000 3.765000 0.455000 ;
      RECT 3.150000  1.525000 3.535000 1.695000 ;
      RECT 3.255000  0.795000 3.425000 1.375000 ;
      RECT 3.255000  1.375000 3.535000 1.525000 ;
      RECT 3.595000  0.455000 3.765000 1.035000 ;
      RECT 3.595000  1.035000 3.875000 1.205000 ;
      RECT 3.685000  2.235000 4.015000 2.635000 ;
      RECT 3.705000  1.205000 3.875000 1.895000 ;
      RECT 3.935000  0.085000 4.105000 0.865000 ;
      RECT 4.105000  1.445000 4.525000 1.715000 ;
      RECT 4.285000  0.415000 4.525000 1.445000 ;
      RECT 4.350000  2.065000 4.520000 2.275000 ;
      RECT 4.350000  2.275000 7.445000 2.445000 ;
      RECT 4.705000  0.265000 5.115000 0.485000 ;
      RECT 4.705000  0.485000 4.915000 0.595000 ;
      RECT 4.705000  0.595000 4.875000 2.105000 ;
      RECT 5.045000  0.720000 5.455000 0.825000 ;
      RECT 5.045000  0.825000 5.255000 0.890000 ;
      RECT 5.045000  0.890000 5.215000 2.275000 ;
      RECT 5.085000  0.655000 5.455000 0.720000 ;
      RECT 5.285000  0.320000 5.455000 0.655000 ;
      RECT 5.395000  1.445000 6.175000 1.615000 ;
      RECT 5.395000  1.615000 5.810000 2.045000 ;
      RECT 5.410000  0.995000 5.835000 1.270000 ;
      RECT 5.625000  0.630000 5.835000 0.995000 ;
      RECT 6.005000  0.255000 7.150000 0.425000 ;
      RECT 6.005000  0.425000 6.175000 1.445000 ;
      RECT 6.345000  0.595000 6.515000 1.935000 ;
      RECT 6.345000  1.935000 8.655000 2.105000 ;
      RECT 6.685000  0.425000 7.150000 0.465000 ;
      RECT 7.025000  0.730000 7.230000 0.945000 ;
      RECT 7.025000  0.945000 7.335000 1.275000 ;
      RECT 7.435000  1.495000 8.255000 1.705000 ;
      RECT 7.475000  0.295000 7.765000 0.735000 ;
      RECT 7.475000  0.735000 8.255000 0.750000 ;
      RECT 7.515000  0.750000 8.255000 0.905000 ;
      RECT 7.855000  2.275000 8.190000 2.635000 ;
      RECT 7.935000  0.085000 8.105000 0.565000 ;
      RECT 8.085000  0.905000 8.255000 0.995000 ;
      RECT 8.085000  0.995000 8.315000 1.325000 ;
      RECT 8.085000  1.325000 8.255000 1.495000 ;
      RECT 8.170000  1.875000 8.655000 1.935000 ;
      RECT 8.355000  0.255000 8.655000 0.585000 ;
      RECT 8.360000  2.105000 8.655000 2.465000 ;
      RECT 8.485000  0.585000 8.655000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  1.445000 3.535000 1.615000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  0.765000 4.455000 0.935000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  0.425000 4.915000 0.595000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  0.765000 5.835000 0.935000 ;
      RECT 5.665000  1.445000 5.835000 1.615000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  0.765000 7.215000 0.935000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  0.425000 7.675000 0.595000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
    LAYER met1 ;
      RECT 3.305000 1.415000 3.595000 1.460000 ;
      RECT 3.305000 1.460000 5.895000 1.600000 ;
      RECT 3.305000 1.600000 3.595000 1.645000 ;
      RECT 4.225000 0.735000 4.515000 0.780000 ;
      RECT 4.225000 0.780000 7.275000 0.920000 ;
      RECT 4.225000 0.920000 4.515000 0.965000 ;
      RECT 4.685000 0.395000 4.975000 0.440000 ;
      RECT 4.685000 0.440000 7.735000 0.580000 ;
      RECT 4.685000 0.580000 4.975000 0.625000 ;
      RECT 5.605000 0.735000 5.895000 0.780000 ;
      RECT 5.605000 0.920000 5.895000 0.965000 ;
      RECT 5.605000 1.415000 5.895000 1.460000 ;
      RECT 5.605000 1.600000 5.895000 1.645000 ;
      RECT 6.985000 0.735000 7.275000 0.780000 ;
      RECT 6.985000 0.920000 7.275000 0.965000 ;
      RECT 7.445000 0.395000 7.735000 0.440000 ;
      RECT 7.445000 0.580000 7.735000 0.625000 ;
  END
END sky130_fd_sc_hd__xnor3_2
MACRO sky130_fd_sc_hd__xnor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.425000 1.075000 8.835000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.605000 0.995000 7.775000 1.445000 ;
        RECT 7.605000 1.445000 8.185000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.995000 1.075000 3.560000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.375000 0.875000 0.995000 ;
        RECT 0.625000 0.995000 1.710000 1.325000 ;
        RECT 0.625000 1.325000 0.955000 2.425000 ;
        RECT 1.465000 0.350000 1.725000 0.925000 ;
        RECT 1.465000 0.925000 1.710000 0.995000 ;
        RECT 1.465000 1.325000 1.710000 1.440000 ;
        RECT 1.465000 1.440000 1.745000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.285000  0.085000 0.455000 0.735000 ;
      RECT 0.285000  1.490000 0.455000 2.635000 ;
      RECT 1.125000  0.085000 1.295000 0.735000 ;
      RECT 1.125000  1.495000 1.295000 2.635000 ;
      RECT 1.880000  0.995000 2.085000 1.325000 ;
      RECT 1.895000  0.085000 2.145000 0.525000 ;
      RECT 1.910000  0.695000 2.485000 0.865000 ;
      RECT 1.910000  0.865000 2.085000 0.995000 ;
      RECT 1.915000  1.325000 2.085000 1.875000 ;
      RECT 1.915000  1.875000 2.600000 2.045000 ;
      RECT 1.915000  2.215000 2.250000 2.635000 ;
      RECT 2.315000  0.255000 3.885000 0.425000 ;
      RECT 2.315000  0.425000 2.485000 0.695000 ;
      RECT 2.315000  1.535000 3.900000 1.705000 ;
      RECT 2.430000  2.045000 2.600000 2.235000 ;
      RECT 2.430000  2.235000 3.900000 2.405000 ;
      RECT 2.655000  0.595000 2.825000 1.535000 ;
      RECT 2.940000  1.895000 5.440000 2.065000 ;
      RECT 3.125000  0.625000 4.345000 0.795000 ;
      RECT 3.125000  0.795000 3.505000 0.905000 ;
      RECT 3.450000  0.425000 3.885000 0.455000 ;
      RECT 3.730000  0.995000 4.005000 1.325000 ;
      RECT 3.730000  1.325000 3.900000 1.535000 ;
      RECT 4.055000  0.285000 4.685000 0.455000 ;
      RECT 4.070000  1.525000 4.455000 1.695000 ;
      RECT 4.175000  0.795000 4.345000 1.375000 ;
      RECT 4.175000  1.375000 4.455000 1.525000 ;
      RECT 4.515000  0.455000 4.685000 1.035000 ;
      RECT 4.515000  1.035000 4.795000 1.205000 ;
      RECT 4.605000  2.235000 4.935000 2.635000 ;
      RECT 4.625000  1.205000 4.795000 1.895000 ;
      RECT 4.855000  0.085000 5.025000 0.865000 ;
      RECT 5.025000  1.445000 5.445000 1.715000 ;
      RECT 5.205000  0.415000 5.445000 1.445000 ;
      RECT 5.270000  2.065000 5.440000 2.275000 ;
      RECT 5.270000  2.275000 8.365000 2.445000 ;
      RECT 5.625000  0.265000 6.035000 0.485000 ;
      RECT 5.625000  0.485000 5.835000 0.595000 ;
      RECT 5.625000  0.595000 5.795000 2.105000 ;
      RECT 5.965000  0.720000 6.375000 0.825000 ;
      RECT 5.965000  0.825000 6.175000 0.890000 ;
      RECT 5.965000  0.890000 6.135000 2.275000 ;
      RECT 6.005000  0.655000 6.375000 0.720000 ;
      RECT 6.205000  0.320000 6.375000 0.655000 ;
      RECT 6.315000  1.445000 7.095000 1.615000 ;
      RECT 6.315000  1.615000 6.730000 2.045000 ;
      RECT 6.330000  0.995000 6.755000 1.270000 ;
      RECT 6.545000  0.630000 6.755000 0.995000 ;
      RECT 6.925000  0.255000 8.070000 0.425000 ;
      RECT 6.925000  0.425000 7.095000 1.445000 ;
      RECT 7.265000  0.595000 7.435000 1.935000 ;
      RECT 7.265000  1.935000 9.575000 2.105000 ;
      RECT 7.605000  0.425000 8.070000 0.465000 ;
      RECT 7.945000  0.730000 8.150000 0.945000 ;
      RECT 7.945000  0.945000 8.255000 1.275000 ;
      RECT 8.355000  1.495000 9.175000 1.705000 ;
      RECT 8.395000  0.295000 8.685000 0.735000 ;
      RECT 8.395000  0.735000 9.175000 0.750000 ;
      RECT 8.435000  0.750000 9.175000 0.905000 ;
      RECT 8.775000  2.275000 9.110000 2.635000 ;
      RECT 8.855000  0.085000 9.025000 0.565000 ;
      RECT 9.005000  0.905000 9.175000 0.995000 ;
      RECT 9.005000  0.995000 9.235000 1.325000 ;
      RECT 9.005000  1.325000 9.175000 1.495000 ;
      RECT 9.090000  1.875000 9.575000 1.935000 ;
      RECT 9.275000  0.255000 9.575000 0.585000 ;
      RECT 9.280000  2.105000 9.575000 2.465000 ;
      RECT 9.405000  0.585000 9.575000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  1.445000 4.455000 1.615000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  0.765000 5.375000 0.935000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  0.425000 5.835000 0.595000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  0.765000 6.755000 0.935000 ;
      RECT 6.585000  1.445000 6.755000 1.615000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  0.765000 8.135000 0.935000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  0.425000 8.595000 0.595000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 4.225000 1.415000 4.515000 1.460000 ;
      RECT 4.225000 1.460000 6.815000 1.600000 ;
      RECT 4.225000 1.600000 4.515000 1.645000 ;
      RECT 5.145000 0.735000 5.435000 0.780000 ;
      RECT 5.145000 0.780000 8.195000 0.920000 ;
      RECT 5.145000 0.920000 5.435000 0.965000 ;
      RECT 5.605000 0.395000 5.895000 0.440000 ;
      RECT 5.605000 0.440000 8.655000 0.580000 ;
      RECT 5.605000 0.580000 5.895000 0.625000 ;
      RECT 6.525000 0.735000 6.815000 0.780000 ;
      RECT 6.525000 0.920000 6.815000 0.965000 ;
      RECT 6.525000 1.415000 6.815000 1.460000 ;
      RECT 6.525000 1.600000 6.815000 1.645000 ;
      RECT 7.905000 0.735000 8.195000 0.780000 ;
      RECT 7.905000 0.920000 8.195000 0.965000 ;
      RECT 8.365000 0.395000 8.655000 0.440000 ;
      RECT 8.365000 0.580000 8.655000 0.625000 ;
  END
END sky130_fd_sc_hd__xnor3_4
MACRO sky130_fd_sc_hd__xnor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.045000 1.075000 7.455000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.225000 0.995000 6.395000 1.445000 ;
        RECT 6.225000 1.445000 6.805000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.615000 1.075000 2.180000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.345000 0.925000 ;
        RECT 0.085000 0.925000 0.330000 1.440000 ;
        RECT 0.085000 1.440000 0.365000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.500000  0.995000 0.705000 1.325000 ;
      RECT 0.515000  0.085000 0.765000 0.525000 ;
      RECT 0.530000  0.695000 1.105000 0.865000 ;
      RECT 0.530000  0.865000 0.705000 0.995000 ;
      RECT 0.535000  1.325000 0.705000 1.875000 ;
      RECT 0.535000  1.875000 1.220000 2.045000 ;
      RECT 0.535000  2.215000 0.870000 2.635000 ;
      RECT 0.935000  0.255000 2.505000 0.425000 ;
      RECT 0.935000  0.425000 1.105000 0.695000 ;
      RECT 0.935000  1.535000 2.520000 1.705000 ;
      RECT 1.050000  2.045000 1.220000 2.235000 ;
      RECT 1.050000  2.235000 2.520000 2.405000 ;
      RECT 1.275000  0.595000 1.445000 1.535000 ;
      RECT 1.560000  1.895000 4.060000 2.065000 ;
      RECT 1.745000  0.625000 2.965000 0.795000 ;
      RECT 1.745000  0.795000 2.125000 0.905000 ;
      RECT 2.070000  0.425000 2.505000 0.455000 ;
      RECT 2.350000  0.995000 2.625000 1.325000 ;
      RECT 2.350000  1.325000 2.520000 1.535000 ;
      RECT 2.675000  0.285000 3.305000 0.455000 ;
      RECT 2.690000  1.525000 3.075000 1.695000 ;
      RECT 2.795000  0.795000 2.965000 1.375000 ;
      RECT 2.795000  1.375000 3.075000 1.525000 ;
      RECT 3.135000  0.455000 3.305000 1.035000 ;
      RECT 3.135000  1.035000 3.415000 1.205000 ;
      RECT 3.225000  2.235000 3.555000 2.635000 ;
      RECT 3.245000  1.205000 3.415000 1.895000 ;
      RECT 3.475000  0.085000 3.645000 0.865000 ;
      RECT 3.645000  1.445000 4.065000 1.715000 ;
      RECT 3.825000  0.415000 4.065000 1.445000 ;
      RECT 3.890000  2.065000 4.060000 2.275000 ;
      RECT 3.890000  2.275000 6.985000 2.445000 ;
      RECT 4.245000  0.265000 4.655000 0.485000 ;
      RECT 4.245000  0.485000 4.455000 0.595000 ;
      RECT 4.245000  0.595000 4.415000 2.105000 ;
      RECT 4.585000  0.720000 4.995000 0.825000 ;
      RECT 4.585000  0.825000 4.795000 0.890000 ;
      RECT 4.585000  0.890000 4.755000 2.275000 ;
      RECT 4.625000  0.655000 4.995000 0.720000 ;
      RECT 4.825000  0.320000 4.995000 0.655000 ;
      RECT 4.935000  1.445000 5.715000 1.615000 ;
      RECT 4.935000  1.615000 5.350000 2.045000 ;
      RECT 4.950000  0.995000 5.375000 1.270000 ;
      RECT 5.165000  0.630000 5.375000 0.995000 ;
      RECT 5.545000  0.255000 6.690000 0.425000 ;
      RECT 5.545000  0.425000 5.715000 1.445000 ;
      RECT 5.885000  0.595000 6.055000 1.935000 ;
      RECT 5.885000  1.935000 8.195000 2.105000 ;
      RECT 6.225000  0.425000 6.690000 0.465000 ;
      RECT 6.565000  0.730000 6.770000 0.945000 ;
      RECT 6.565000  0.945000 6.875000 1.275000 ;
      RECT 6.975000  1.495000 7.795000 1.705000 ;
      RECT 7.015000  0.295000 7.305000 0.735000 ;
      RECT 7.015000  0.735000 7.795000 0.750000 ;
      RECT 7.055000  0.750000 7.795000 0.905000 ;
      RECT 7.395000  2.275000 7.730000 2.635000 ;
      RECT 7.475000  0.085000 7.645000 0.565000 ;
      RECT 7.625000  0.905000 7.795000 0.995000 ;
      RECT 7.625000  0.995000 7.855000 1.325000 ;
      RECT 7.625000  1.325000 7.795000 1.495000 ;
      RECT 7.710000  1.875000 8.195000 1.935000 ;
      RECT 7.895000  0.255000 8.195000 0.585000 ;
      RECT 7.900000  2.105000 8.195000 2.465000 ;
      RECT 8.025000  0.585000 8.195000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  1.445000 3.075000 1.615000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  0.765000 3.995000 0.935000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  0.425000 4.455000 0.595000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  0.765000 5.375000 0.935000 ;
      RECT 5.205000  1.445000 5.375000 1.615000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  0.765000 6.755000 0.935000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  0.425000 7.215000 0.595000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 2.845000 1.415000 3.135000 1.460000 ;
      RECT 2.845000 1.460000 5.435000 1.600000 ;
      RECT 2.845000 1.600000 3.135000 1.645000 ;
      RECT 3.765000 0.735000 4.055000 0.780000 ;
      RECT 3.765000 0.780000 6.815000 0.920000 ;
      RECT 3.765000 0.920000 4.055000 0.965000 ;
      RECT 4.225000 0.395000 4.515000 0.440000 ;
      RECT 4.225000 0.440000 7.275000 0.580000 ;
      RECT 4.225000 0.580000 4.515000 0.625000 ;
      RECT 5.145000 0.735000 5.435000 0.780000 ;
      RECT 5.145000 0.920000 5.435000 0.965000 ;
      RECT 5.145000 1.415000 5.435000 1.460000 ;
      RECT 5.145000 1.600000 5.435000 1.645000 ;
      RECT 6.525000 0.735000 6.815000 0.780000 ;
      RECT 6.525000 0.920000 6.815000 0.965000 ;
      RECT 6.985000 0.395000 7.275000 0.440000 ;
      RECT 6.985000 0.580000 7.275000 0.625000 ;
  END
END sky130_fd_sc_hd__xnor3_1
MACRO sky130_fd_sc_hd__o41ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.500000 1.075000 3.080000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.415000 2.330000 2.355000 ;
        RECT 2.000000 1.075000 2.330000 1.415000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 1.075000 1.830000 1.245000 ;
        RECT 1.500000 1.245000 1.820000 2.355000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.990000 1.075000 1.320000 1.245000 ;
        RECT 1.015000 1.245000 1.320000 2.355000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 0.440000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 0.735000 ;
        RECT 0.085000 0.735000 0.780000 0.905000 ;
        RECT 0.515000 1.485000 0.845000 2.465000 ;
        RECT 0.610000 0.905000 0.780000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.445000 0.345000 2.635000 ;
      RECT 0.790000  0.255000 1.120000 0.565000 ;
      RECT 0.950000  0.565000 1.120000 0.735000 ;
      RECT 0.950000  0.735000 2.960000 0.905000 ;
      RECT 1.290000  0.085000 1.540000 0.565000 ;
      RECT 1.710000  0.255000 2.040000 0.735000 ;
      RECT 2.210000  0.085000 2.460000 0.565000 ;
      RECT 2.630000  0.255000 2.960000 0.735000 ;
      RECT 2.630000  1.495000 2.960000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o41ai_1
MACRO sky130_fd_sc_hd__o41ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.155000 1.075000 10.035000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.170000 1.075000 7.940000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.310000 1.075000 5.980000 1.275000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.350000 1.075000 4.020000 1.275000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 1.700000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 2.160000 0.905000 ;
        RECT 0.515000 1.445000 3.885000 1.615000 ;
        RECT 0.515000 1.615000 0.845000 2.465000 ;
        RECT 1.355000 1.615000 1.685000 2.465000 ;
        RECT 1.870000 0.905000 2.160000 1.445000 ;
        RECT 2.715000 1.615000 3.045000 2.125000 ;
        RECT 3.555000 1.615000 3.885000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.255000  2.625000 0.465000 ;
      RECT 0.085000  0.465000  0.345000 0.905000 ;
      RECT 0.085000  1.445000  0.345000 2.635000 ;
      RECT 1.015000  1.835000  1.185000 2.635000 ;
      RECT 1.855000  1.835000  2.105000 2.635000 ;
      RECT 2.295000  1.785000  2.545000 2.295000 ;
      RECT 2.295000  2.295000  4.225000 2.465000 ;
      RECT 2.350000  0.465000  2.625000 0.735000 ;
      RECT 2.350000  0.735000  9.865000 0.905000 ;
      RECT 2.795000  0.085000  2.965000 0.545000 ;
      RECT 3.135000  0.255000  3.465000 0.735000 ;
      RECT 3.215000  1.785000  3.385000 2.295000 ;
      RECT 3.635000  0.085000  3.805000 0.545000 ;
      RECT 3.975000  0.255000  4.305000 0.735000 ;
      RECT 4.055000  1.445000  5.985000 1.615000 ;
      RECT 4.055000  1.615000  4.225000 2.295000 ;
      RECT 4.395000  1.785000  4.645000 2.295000 ;
      RECT 4.395000  2.295000  7.685000 2.465000 ;
      RECT 4.475000  0.085000  4.645000 0.545000 ;
      RECT 4.815000  0.255000  5.145000 0.735000 ;
      RECT 4.815000  1.615000  5.145000 2.125000 ;
      RECT 5.315000  0.085000  5.485000 0.545000 ;
      RECT 5.315000  1.785000  5.485000 2.295000 ;
      RECT 5.655000  0.255000  5.985000 0.735000 ;
      RECT 5.655000  1.615000  5.985000 2.125000 ;
      RECT 6.175000  0.260000  6.505000 0.735000 ;
      RECT 6.175000  1.445000  9.865000 1.615000 ;
      RECT 6.175000  1.615000  6.505000 2.125000 ;
      RECT 6.675000  0.085000  6.845000 0.545000 ;
      RECT 6.675000  1.785000  6.845000 2.295000 ;
      RECT 7.015000  0.260000  7.345000 0.735000 ;
      RECT 7.015000  1.615000  7.345000 2.125000 ;
      RECT 7.515000  0.085000  7.685000 0.545000 ;
      RECT 7.515000  1.785000  7.685000 2.295000 ;
      RECT 7.855000  0.260000  8.185000 0.735000 ;
      RECT 7.855000  1.615000  8.185000 2.465000 ;
      RECT 8.355000  0.085000  8.525000 0.545000 ;
      RECT 8.355000  1.835000  8.525000 2.635000 ;
      RECT 8.695000  0.260000  9.025000 0.735000 ;
      RECT 8.695000  1.615000  9.025000 2.465000 ;
      RECT 9.195000  0.085000  9.365000 0.545000 ;
      RECT 9.195000  1.835000  9.365000 2.635000 ;
      RECT 9.535000  0.260000  9.865000 0.735000 ;
      RECT 9.535000  1.615000  9.865000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__o41ai_4
MACRO sky130_fd_sc_hd__o41ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.720000 1.075000 5.895000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.780000 1.075000 4.540000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.595000 1.075000 3.580000 1.275000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 1.075000 2.325000 1.275000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.075000 0.440000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 0.845000 0.885000 ;
        RECT 0.515000 1.505000 2.205000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 0.610000 0.885000 0.845000 1.445000 ;
        RECT 0.610000 1.445000 2.205000 1.505000 ;
        RECT 1.875000 1.665000 2.205000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.255000 1.265000 0.465000 ;
      RECT 0.085000  0.465000 0.345000 0.905000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 1.015000  0.465000 1.265000 0.735000 ;
      RECT 1.015000  0.735000 5.705000 0.905000 ;
      RECT 1.015000  1.835000 1.265000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.455000  1.835000 1.705000 2.295000 ;
      RECT 1.455000  2.295000 2.545000 2.465000 ;
      RECT 1.875000  0.255000 2.205000 0.735000 ;
      RECT 2.375000  0.085000 2.545000 0.545000 ;
      RECT 2.375000  1.445000 3.465000 1.615000 ;
      RECT 2.375000  1.615000 2.545000 2.295000 ;
      RECT 2.715000  0.255000 3.045000 0.735000 ;
      RECT 2.715000  1.835000 3.045000 2.295000 ;
      RECT 2.715000  2.295000 4.445000 2.465000 ;
      RECT 3.215000  0.085000 3.450000 0.545000 ;
      RECT 3.215000  1.615000 3.465000 2.125000 ;
      RECT 3.695000  0.255000 4.025000 0.735000 ;
      RECT 3.695000  1.445000 5.705000 1.615000 ;
      RECT 3.695000  1.615000 3.945000 2.125000 ;
      RECT 4.115000  1.835000 4.445000 2.295000 ;
      RECT 4.195000  0.085000 4.365000 0.545000 ;
      RECT 4.535000  0.255000 4.865000 0.735000 ;
      RECT 4.615000  1.615000 4.785000 2.465000 ;
      RECT 4.955000  1.785000 5.285000 2.635000 ;
      RECT 5.035000  0.085000 5.205000 0.545000 ;
      RECT 5.375000  0.255000 5.705000 0.735000 ;
      RECT 5.455000  1.615000 5.705000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__o41ai_2
MACRO sky130_fd_sc_hd__o41a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 1.075000 4.515000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.325000 1.075000 3.655000 2.335000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.825000 1.075000 3.155000 2.340000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 1.075000 2.655000 2.340000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775000 1.075000 2.155000 1.325000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.845000 0.880000 ;
        RECT 0.515000 0.880000 0.790000 1.495000 ;
        RECT 0.515000 1.495000 0.845000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.885000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.960000  1.075000 1.600000 1.325000 ;
      RECT 1.015000  0.085000 1.260000 0.885000 ;
      RECT 1.015000  1.495000 1.185000 1.835000 ;
      RECT 1.015000  1.835000 1.525000 2.635000 ;
      RECT 1.355000  1.325000 1.600000 1.495000 ;
      RECT 1.355000  1.495000 2.145000 1.665000 ;
      RECT 1.430000  0.255000 1.785000 0.850000 ;
      RECT 1.430000  0.850000 1.600000 1.075000 ;
      RECT 1.695000  1.665000 2.145000 2.465000 ;
      RECT 1.985000  0.255000 2.315000 0.715000 ;
      RECT 1.985000  0.715000 4.395000 0.905000 ;
      RECT 2.485000  0.085000 2.750000 0.545000 ;
      RECT 2.955000  0.255000 3.285000 0.715000 ;
      RECT 3.505000  0.085000 3.775000 0.545000 ;
      RECT 4.065000  0.255000 4.395000 0.715000 ;
      RECT 4.065000  1.495000 4.395000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__o41a_2
MACRO sky130_fd_sc_hd__o41a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.650000 1.075000 7.735000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.150000 1.075000 6.360000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.330000 1.075000 4.960000 1.275000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.410000 1.075000 4.040000 1.275000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.835000 1.075000 3.165000 1.275000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 1.685000 0.905000 ;
        RECT 0.085000 0.905000 0.345000 1.465000 ;
        RECT 0.085000 1.465000 1.685000 1.665000 ;
        RECT 0.515000 0.255000 0.845000 0.715000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 0.255000 1.685000 0.715000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.545000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  1.075000 2.665000 1.245000 ;
      RECT 0.515000  1.245000 2.545000 1.295000 ;
      RECT 1.015000  0.085000 1.185000 0.545000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.855000  0.085000 2.105000 0.885000 ;
      RECT 1.855000  1.465000 2.025000 2.635000 ;
      RECT 2.195000  1.295000 2.545000 1.445000 ;
      RECT 2.195000  1.445000 3.825000 1.615000 ;
      RECT 2.195000  1.615000 2.545000 2.465000 ;
      RECT 2.295000  0.255000 3.485000 0.465000 ;
      RECT 2.295000  0.635000 3.045000 0.905000 ;
      RECT 2.295000  0.905000 2.665000 1.075000 ;
      RECT 2.715000  1.835000 2.965000 2.635000 ;
      RECT 3.135000  1.835000 3.405000 2.295000 ;
      RECT 3.135000  2.295000 4.325000 2.465000 ;
      RECT 3.235000  0.465000 3.485000 0.735000 ;
      RECT 3.235000  0.735000 7.595000 0.905000 ;
      RECT 3.575000  1.615000 3.825000 2.125000 ;
      RECT 3.655000  0.085000 3.875000 0.545000 ;
      RECT 3.995000  1.445000 5.165000 1.615000 ;
      RECT 3.995000  1.615000 4.325000 2.295000 ;
      RECT 4.075000  0.255000 4.245000 0.735000 ;
      RECT 4.445000  0.085000 4.715000 0.545000 ;
      RECT 4.495000  1.785000 4.665000 2.295000 ;
      RECT 4.495000  2.295000 6.145000 2.465000 ;
      RECT 4.835000  1.615000 5.165000 2.115000 ;
      RECT 4.915000  0.255000 5.085000 0.735000 ;
      RECT 5.305000  0.085000 5.915000 0.545000 ;
      RECT 5.395000  1.445000 7.595000 1.615000 ;
      RECT 5.395000  1.615000 5.645000 2.115000 ;
      RECT 5.815000  1.785000 6.145000 2.295000 ;
      RECT 6.240000  0.255000 6.410000 0.735000 ;
      RECT 6.315000  1.615000 6.485000 2.455000 ;
      RECT 6.655000  1.785000 6.985000 2.635000 ;
      RECT 6.685000  0.085000 6.955000 0.545000 ;
      RECT 7.265000  0.255000 7.595000 0.735000 ;
      RECT 7.265000  1.615000 7.595000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__o41a_4
MACRO sky130_fd_sc_hd__o41a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.075000 3.995000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.075000 3.275000 2.390000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.075000 2.735000 2.390000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.865000 1.075000 2.195000 2.390000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275000 1.075000 1.695000 1.285000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.672000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 0.885000 ;
        RECT 0.085000 0.885000 0.355000 1.455000 ;
        RECT 0.085000 1.455000 0.610000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.525000  1.075000 1.105000 1.285000 ;
      RECT 0.715000  0.085000 0.885000 0.545000 ;
      RECT 0.735000  0.715000 1.485000 0.905000 ;
      RECT 0.735000  0.905000 1.105000 1.075000 ;
      RECT 0.845000  1.285000 1.105000 1.455000 ;
      RECT 0.845000  1.455000 1.595000 1.745000 ;
      RECT 0.845000  1.915000 1.175000 2.635000 ;
      RECT 1.155000  0.270000 1.485000 0.715000 ;
      RECT 1.345000  1.745000 1.595000 2.465000 ;
      RECT 1.655000  0.415000 1.825000 0.735000 ;
      RECT 1.655000  0.735000 3.955000 0.905000 ;
      RECT 2.050000  0.085000 2.380000 0.545000 ;
      RECT 2.580000  0.255000 2.910000 0.735000 ;
      RECT 3.125000  0.085000 3.455000 0.545000 ;
      RECT 3.605000  1.515000 3.935000 2.635000 ;
      RECT 3.625000  0.255000 3.955000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o41a_1
MACRO sky130_fd_sc_hd__dlxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 0.955000 1.685000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.140000 0.255000 5.490000 0.820000 ;
        RECT 5.140000 1.670000 5.490000 2.455000 ;
        RECT 5.320000 0.820000 5.490000 1.670000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.555000 0.255000 6.815000 0.825000 ;
        RECT 6.555000 1.445000 6.815000 2.465000 ;
        RECT 6.600000 0.825000 6.815000 1.445000 ;
    END
  END Q_N
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.430000  1.495000 2.115000 1.665000 ;
      RECT 1.430000  1.665000 1.795000 2.415000 ;
      RECT 1.510000  0.345000 1.705000 0.615000 ;
      RECT 1.510000  0.615000 2.135000 0.785000 ;
      RECT 1.855000  0.785000 2.135000 0.875000 ;
      RECT 1.855000  0.875000 2.335000 1.235000 ;
      RECT 1.855000  1.235000 2.115000 1.495000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.965000  1.835000 2.245000 2.635000 ;
      RECT 2.465000  1.355000 2.795000 1.685000 ;
      RECT 2.580000  0.705000 3.135000 1.065000 ;
      RECT 2.750000  2.255000 3.610000 2.425000 ;
      RECT 2.800000  0.365000 3.475000 0.535000 ;
      RECT 2.965000  1.065000 3.135000 1.575000 ;
      RECT 2.965000  1.575000 3.290000 1.910000 ;
      RECT 2.965000  1.910000 3.195000 1.995000 ;
      RECT 3.305000  0.535000 3.475000 0.995000 ;
      RECT 3.305000  0.995000 4.175000 1.165000 ;
      RECT 3.425000  2.035000 3.650000 2.065000 ;
      RECT 3.425000  2.065000 3.630000 2.090000 ;
      RECT 3.425000  2.090000 3.610000 2.255000 ;
      RECT 3.430000  2.020000 3.650000 2.035000 ;
      RECT 3.435000  2.010000 3.650000 2.020000 ;
      RECT 3.440000  1.995000 3.650000 2.010000 ;
      RECT 3.460000  1.165000 4.175000 1.325000 ;
      RECT 3.460000  1.325000 3.650000 1.995000 ;
      RECT 3.700000  0.085000 4.045000 0.530000 ;
      RECT 3.780000  2.175000 3.980000 2.635000 ;
      RECT 3.820000  1.535000 4.515000 1.865000 ;
      RECT 4.285000  0.415000 4.550000 0.745000 ;
      RECT 4.285000  1.865000 4.515000 2.435000 ;
      RECT 4.345000  0.745000 4.550000 0.995000 ;
      RECT 4.345000  0.995000 5.150000 1.325000 ;
      RECT 4.345000  1.325000 4.515000 1.535000 ;
      RECT 4.685000  1.570000 4.970000 2.635000 ;
      RECT 4.720000  0.085000 4.970000 0.715000 ;
      RECT 5.660000  0.255000 5.910000 0.995000 ;
      RECT 5.660000  0.995000 6.430000 1.325000 ;
      RECT 5.660000  1.325000 5.910000 2.465000 ;
      RECT 6.090000  0.085000 6.385000 0.545000 ;
      RECT 6.090000  1.835000 6.385000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.555000  1.445000 2.725000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.965000  1.785000 3.135000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 2.785000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 3.195000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.495000 1.415000 2.785000 1.460000 ;
      RECT 2.495000 1.600000 2.785000 1.645000 ;
      RECT 2.905000 1.755000 3.195000 1.800000 ;
      RECT 2.905000 1.940000 3.195000 1.985000 ;
  END
END sky130_fd_sc_hd__dlxbp_1
MACRO sky130_fd_sc_hd__o211ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505000 1.075000 4.455000 1.245000 ;
        RECT 3.560000 1.245000 4.455000 1.295000 ;
        RECT 4.115000 0.765000 4.455000 1.075000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365000 1.075000 3.335000 1.355000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.075000 1.905000 1.365000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.375000 1.970000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.022000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.670000 0.875000 1.540000 ;
        RECT 0.545000 1.540000 3.155000 1.710000 ;
        RECT 0.545000 1.710000 0.805000 2.465000 ;
        RECT 1.475000 1.710000 1.665000 2.465000 ;
        RECT 2.825000 1.710000 3.155000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.095000  0.255000 2.165000 0.445000 ;
      RECT 0.115000  2.175000 0.375000 2.635000 ;
      RECT 0.975000  1.915000 1.305000 2.635000 ;
      RECT 1.045000  0.445000 2.165000 0.465000 ;
      RECT 1.045000  0.465000 1.235000 0.890000 ;
      RECT 1.405000  0.635000 3.945000 0.845000 ;
      RECT 1.835000  1.915000 2.165000 2.635000 ;
      RECT 2.395000  0.085000 2.725000 0.445000 ;
      RECT 2.395000  2.100000 2.655000 2.295000 ;
      RECT 2.395000  2.295000 3.515000 2.465000 ;
      RECT 3.255000  0.085000 3.585000 0.445000 ;
      RECT 3.325000  1.525000 4.445000 1.695000 ;
      RECT 3.325000  1.695000 3.515000 2.295000 ;
      RECT 3.685000  1.865000 4.015000 2.635000 ;
      RECT 3.755000  0.515000 3.945000 0.635000 ;
      RECT 4.115000  0.085000 4.445000 0.445000 ;
      RECT 4.185000  1.695000 4.445000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__o211ai_2
MACRO sky130_fd_sc_hd__o211ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.395000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.995000 0.980000 1.325000 ;
        RECT 0.605000 1.325000 0.775000 2.250000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.300000 0.995000 1.795000 1.325000 ;
        RECT 1.470000 1.325000 1.795000 1.615000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 1.075000 2.300000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.418250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 1.595000 1.275000 1.815000 ;
        RECT 0.945000 1.815000 2.675000 2.045000 ;
        RECT 0.945000 2.045000 1.275000 2.445000 ;
        RECT 1.965000 0.255000 2.675000 0.845000 ;
        RECT 1.975000 2.045000 2.675000 2.465000 ;
        RECT 2.470000 0.845000 2.675000 1.815000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  0.255000 0.425000 0.615000 ;
      RECT 0.095000  0.615000 1.455000 0.825000 ;
      RECT 0.095000  1.575000 0.425000 2.635000 ;
      RECT 0.595000  0.085000 0.925000 0.445000 ;
      RECT 1.125000  0.255000 1.455000 0.615000 ;
      RECT 1.445000  2.275000 1.775000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__o211ai_1
MACRO sky130_fd_sc_hd__o211ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.400000 1.075000 1.410000 1.330000 ;
        RECT 0.965000 1.330000 1.410000 1.515000 ;
        RECT 0.965000 1.515000 3.630000 1.685000 ;
        RECT 3.350000 0.995000 3.630000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.705000 1.075000 3.180000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.800000 0.995000 4.975000 1.410000 ;
        RECT 4.260000 1.410000 4.975000 1.515000 ;
        RECT 4.260000 1.515000 7.000000 1.685000 ;
        RECT 6.830000 0.995000 7.000000 1.515000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.370000 1.075000 6.440000 1.345000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.001000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 1.855000 7.680000 2.025000 ;
        RECT 1.805000 2.025000 3.470000 2.105000 ;
        RECT 4.045000 2.025000 7.680000 2.105000 ;
        RECT 5.280000 0.270000 6.735000 0.450000 ;
        RECT 6.565000 0.450000 6.735000 0.655000 ;
        RECT 6.565000 0.655000 7.350000 0.825000 ;
        RECT 7.170000 0.825000 7.350000 1.340000 ;
        RECT 7.170000 1.340000 7.680000 1.855000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.090000  1.665000 0.385000 2.635000 ;
      RECT 0.155000  0.535000 0.355000 0.625000 ;
      RECT 0.155000  0.625000 1.240000 0.695000 ;
      RECT 0.155000  0.695000 3.835000 0.795000 ;
      RECT 0.155000  0.795000 3.130000 0.865000 ;
      RECT 0.155000  0.865000 1.795000 0.905000 ;
      RECT 0.525000  0.085000 0.855000 0.445000 ;
      RECT 0.555000  1.860000 0.775000 1.935000 ;
      RECT 0.555000  1.935000 1.635000 2.105000 ;
      RECT 0.555000  2.105000 0.775000 2.190000 ;
      RECT 0.955000  2.275000 1.285000 2.635000 ;
      RECT 1.025000  0.425000 1.240000 0.625000 ;
      RECT 1.455000  2.105000 1.635000 2.275000 ;
      RECT 1.455000  2.275000 3.435000 2.465000 ;
      RECT 1.465000  0.085000 1.635000 0.525000 ;
      RECT 1.775000  0.625000 3.835000 0.695000 ;
      RECT 2.245000  0.085000 2.575000 0.445000 ;
      RECT 3.105000  0.085000 3.435000 0.445000 ;
      RECT 3.605000  0.255000 4.920000 0.455000 ;
      RECT 3.605000  0.455000 3.835000 0.625000 ;
      RECT 3.615000  2.195000 3.885000 2.635000 ;
      RECT 4.005000  0.635000 6.170000 0.815000 ;
      RECT 4.435000  2.275000 4.765000 2.635000 ;
      RECT 5.280000  2.275000 5.610000 2.635000 ;
      RECT 6.120000  2.275000 6.455000 2.635000 ;
      RECT 6.980000  0.310000 7.680000 0.480000 ;
      RECT 7.355000  2.275000 7.685000 2.635000 ;
      RECT 7.510000  0.480000 7.680000 0.595000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  0.425000 1.240000 0.595000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.510000  0.425000 7.680000 0.595000 ;
    LAYER met1 ;
      RECT 1.010000 0.395000 1.300000 0.440000 ;
      RECT 1.010000 0.440000 7.740000 0.580000 ;
      RECT 1.010000 0.580000 1.300000 0.625000 ;
      RECT 7.450000 0.395000 7.740000 0.440000 ;
      RECT 7.450000 0.580000 7.740000 0.625000 ;
  END
END sky130_fd_sc_hd__o211ai_4
MACRO sky130_fd_sc_hd__dfbbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfbbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.750000 1.005000 2.160000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.615000 0.255000 11.875000 0.825000 ;
        RECT 11.615000 1.445000 11.875000 2.465000 ;
        RECT 11.660000 0.825000 11.875000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.200000 0.255000 10.485000 0.715000 ;
        RECT 10.200000 1.630000 10.485000 2.465000 ;
        RECT 10.280000 0.715000 10.485000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.315000 1.095000 9.690000 1.325000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.590000 0.735000 4.000000 0.965000 ;
        RECT 3.590000 0.965000 3.920000 1.065000 ;
      LAYER mcon ;
        RECT 3.830000 0.765000 4.000000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.460000 0.735000 7.835000 1.065000 ;
      LAYER mcon ;
        RECT 7.510000 0.765000 7.680000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.770000 0.735000 4.060000 0.780000 ;
        RECT 3.770000 0.780000 7.740000 0.920000 ;
        RECT 3.770000 0.920000 4.060000 0.965000 ;
        RECT 7.450000 0.735000 7.740000 0.780000 ;
        RECT 7.450000 0.920000 7.740000 0.965000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.085000  0.345000  0.345000 0.635000 ;
      RECT  0.085000  0.635000  0.840000 0.805000 ;
      RECT  0.085000  1.795000  0.840000 1.965000 ;
      RECT  0.085000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.240000 2.465000 ;
      RECT  1.410000  0.635000  2.125000 0.825000 ;
      RECT  1.410000  0.825000  1.580000 1.795000 ;
      RECT  1.410000  1.795000  2.125000 1.965000 ;
      RECT  1.435000  0.085000  1.785000 0.465000 ;
      RECT  1.435000  2.135000  1.785000 2.635000 ;
      RECT  1.955000  0.305000  2.125000 0.635000 ;
      RECT  1.955000  1.965000  2.125000 2.465000 ;
      RECT  2.330000  0.705000  2.550000 1.575000 ;
      RECT  2.330000  1.575000  2.830000 1.955000 ;
      RECT  2.340000  2.250000  3.170000 2.420000 ;
      RECT  2.405000  0.265000  3.400000 0.465000 ;
      RECT  2.730000  0.645000  3.060000 1.015000 ;
      RECT  3.000000  1.195000  3.400000 1.235000 ;
      RECT  3.000000  1.235000  4.350000 1.405000 ;
      RECT  3.000000  1.405000  3.170000 2.250000 ;
      RECT  3.230000  0.465000  3.400000 1.195000 ;
      RECT  3.340000  1.575000  3.590000 1.785000 ;
      RECT  3.340000  1.785000  4.690000 2.035000 ;
      RECT  3.410000  2.205000  3.790000 2.635000 ;
      RECT  3.570000  0.085000  3.740000 0.525000 ;
      RECT  3.910000  0.255000  5.080000 0.425000 ;
      RECT  3.910000  0.425000  4.240000 0.545000 ;
      RECT  4.090000  2.035000  4.260000 2.375000 ;
      RECT  4.100000  1.405000  4.350000 1.485000 ;
      RECT  4.130000  1.155000  4.350000 1.235000 ;
      RECT  4.410000  0.595000  4.740000 0.765000 ;
      RECT  4.520000  0.765000  4.740000 0.895000 ;
      RECT  4.520000  0.895000  5.830000 1.065000 ;
      RECT  4.520000  1.065000  4.690000 1.785000 ;
      RECT  4.860000  1.235000  5.190000 1.415000 ;
      RECT  4.860000  1.415000  5.865000 1.655000 ;
      RECT  4.880000  1.915000  5.210000 2.635000 ;
      RECT  4.910000  0.425000  5.080000 0.715000 ;
      RECT  5.350000  0.085000  5.680000 0.465000 ;
      RECT  5.500000  1.065000  5.830000 1.235000 ;
      RECT  6.065000  1.575000  6.300000 1.985000 ;
      RECT  6.125000  0.705000  6.410000 1.125000 ;
      RECT  6.125000  1.125000  6.745000 1.305000 ;
      RECT  6.255000  2.250000  7.085000 2.420000 ;
      RECT  6.320000  0.265000  7.085000 0.465000 ;
      RECT  6.540000  1.305000  6.745000 1.905000 ;
      RECT  6.915000  0.465000  7.085000 1.235000 ;
      RECT  6.915000  1.235000  8.265000 1.405000 ;
      RECT  6.915000  1.405000  7.085000 2.250000 ;
      RECT  7.255000  1.575000  7.505000 1.915000 ;
      RECT  7.255000  1.915000 10.030000 2.085000 ;
      RECT  7.265000  0.085000  7.525000 0.525000 ;
      RECT  7.325000  2.255000  7.705000 2.635000 ;
      RECT  7.785000  0.255000  8.955000 0.425000 ;
      RECT  7.785000  0.425000  8.115000 0.545000 ;
      RECT  7.945000  2.085000  8.115000 2.375000 ;
      RECT  8.045000  1.075000  8.265000 1.235000 ;
      RECT  8.285000  0.595000  8.615000 0.780000 ;
      RECT  8.435000  0.780000  8.615000 1.915000 ;
      RECT  8.645000  2.255000 10.030000 2.635000 ;
      RECT  8.785000  0.425000  8.955000 0.585000 ;
      RECT  8.785000  0.755000  9.475000 0.925000 ;
      RECT  8.785000  0.925000  9.060000 1.575000 ;
      RECT  8.785000  1.575000  9.545000 1.745000 ;
      RECT  9.240000  0.265000  9.475000 0.755000 ;
      RECT  9.700000  0.085000 10.030000 0.805000 ;
      RECT  9.860000  0.995000 10.110000 1.325000 ;
      RECT  9.860000  1.325000 10.030000 1.915000 ;
      RECT 10.655000  0.255000 10.970000 0.995000 ;
      RECT 10.655000  0.995000 11.490000 1.325000 ;
      RECT 10.655000  1.325000 10.970000 2.415000 ;
      RECT 11.150000  0.085000 11.445000 0.545000 ;
      RECT 11.150000  1.765000 11.445000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.610000  1.785000  0.780000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.070000  0.765000  1.240000 0.935000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.450000  1.785000  2.620000 1.955000 ;
      RECT  2.890000  0.765000  3.060000 0.935000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.670000  1.445000  5.840000 1.615000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.130000  1.105000  6.300000 1.275000 ;
      RECT  6.130000  1.785000  6.300000 1.955000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.890000  1.445000  9.060000 1.615000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.755000 0.840000 1.800000 ;
      RECT 0.550000 1.800000 6.360000 1.940000 ;
      RECT 0.550000 1.940000 0.840000 1.985000 ;
      RECT 1.010000 0.735000 1.300000 0.780000 ;
      RECT 1.010000 0.780000 3.120000 0.920000 ;
      RECT 1.010000 0.920000 1.300000 0.965000 ;
      RECT 2.390000 1.755000 2.680000 1.800000 ;
      RECT 2.390000 1.940000 2.680000 1.985000 ;
      RECT 2.830000 0.735000 3.120000 0.780000 ;
      RECT 2.830000 0.920000 3.120000 0.965000 ;
      RECT 2.925000 0.965000 3.120000 1.120000 ;
      RECT 2.925000 1.120000 6.360000 1.260000 ;
      RECT 5.610000 1.415000 5.900000 1.460000 ;
      RECT 5.610000 1.460000 9.120000 1.600000 ;
      RECT 5.610000 1.600000 5.900000 1.645000 ;
      RECT 6.070000 1.075000 6.360000 1.120000 ;
      RECT 6.070000 1.260000 6.360000 1.305000 ;
      RECT 6.070000 1.755000 6.360000 1.800000 ;
      RECT 6.070000 1.940000 6.360000 1.985000 ;
      RECT 8.830000 1.415000 9.120000 1.460000 ;
      RECT 8.830000 1.600000 9.120000 1.645000 ;
  END
END sky130_fd_sc_hd__dfbbp_1
MACRO sky130_fd_sc_hd__dlxtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.955000 1.765000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.175000 0.415000 5.435000 0.745000 ;
        RECT 5.175000 1.670000 5.435000 2.455000 ;
        RECT 5.265000 0.745000 5.435000 1.670000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.430000  1.495000 2.115000 1.665000 ;
      RECT 1.430000  1.665000 1.785000 2.415000 ;
      RECT 1.510000  0.345000 1.705000 0.615000 ;
      RECT 1.510000  0.615000 2.115000 0.765000 ;
      RECT 1.510000  0.765000 2.320000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.945000  0.785000 2.320000 1.235000 ;
      RECT 1.945000  1.235000 2.115000 1.495000 ;
      RECT 1.955000  1.835000 2.245000 2.635000 ;
      RECT 2.445000  1.355000 2.780000 2.005000 ;
      RECT 2.560000  0.735000 3.265000 1.040000 ;
      RECT 2.745000  2.255000 3.605000 2.425000 ;
      RECT 2.765000  0.365000 3.605000 0.535000 ;
      RECT 2.950000  1.040000 3.265000 1.560000 ;
      RECT 2.950000  1.560000 3.285000 1.910000 ;
      RECT 3.295000  2.090000 3.620000 2.105000 ;
      RECT 3.295000  2.105000 3.605000 2.255000 ;
      RECT 3.390000  2.045000 3.645000 2.065000 ;
      RECT 3.390000  2.065000 3.630000 2.085000 ;
      RECT 3.390000  2.085000 3.620000 2.090000 ;
      RECT 3.405000  2.035000 3.645000 2.045000 ;
      RECT 3.430000  2.010000 3.645000 2.035000 ;
      RECT 3.435000  0.535000 3.605000 0.995000 ;
      RECT 3.435000  0.995000 4.200000 1.325000 ;
      RECT 3.435000  1.325000 3.645000 1.450000 ;
      RECT 3.455000  1.450000 3.645000 2.010000 ;
      RECT 3.775000  0.085000 4.045000 0.545000 ;
      RECT 3.775000  2.175000 4.095000 2.635000 ;
      RECT 3.815000  1.535000 4.540000 1.865000 ;
      RECT 4.295000  0.260000 4.540000 0.720000 ;
      RECT 4.295000  1.865000 4.540000 2.435000 ;
      RECT 4.370000  0.720000 4.540000 0.995000 ;
      RECT 4.370000  0.995000 5.095000 1.325000 ;
      RECT 4.370000  1.325000 4.540000 1.535000 ;
      RECT 4.720000  1.570000 5.005000 2.635000 ;
      RECT 4.755000  0.085000 4.980000 0.715000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  1.785000 2.615000 1.955000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.950000  1.445000 3.120000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.180000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.675000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.385000 1.755000 2.675000 1.800000 ;
      RECT 2.385000 1.940000 2.675000 1.985000 ;
      RECT 2.890000 1.415000 3.180000 1.460000 ;
      RECT 2.890000 1.600000 3.180000 1.645000 ;
  END
END sky130_fd_sc_hd__dlxtn_1
MACRO sky130_fd_sc_hd__dlxtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 0.955000 1.810000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.215000 0.415000 5.465000 0.685000 ;
        RECT 5.215000 0.685000 5.500000 0.825000 ;
        RECT 5.215000 1.495000 5.500000 1.640000 ;
        RECT 5.215000 1.640000 5.465000 2.455000 ;
        RECT 5.330000 0.825000 5.500000 0.995000 ;
        RECT 5.330000 0.995000 5.895000 1.325000 ;
        RECT 5.330000 1.325000 5.500000 1.495000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.475000  1.495000 2.160000 1.665000 ;
      RECT 1.475000  1.665000 1.805000 2.415000 ;
      RECT 1.555000  0.345000 1.725000 0.615000 ;
      RECT 1.555000  0.615000 2.160000 0.765000 ;
      RECT 1.555000  0.765000 2.360000 0.785000 ;
      RECT 1.895000  0.085000 2.225000 0.445000 ;
      RECT 1.975000  1.835000 2.290000 2.635000 ;
      RECT 1.990000  0.785000 2.360000 1.095000 ;
      RECT 1.990000  1.095000 2.160000 1.495000 ;
      RECT 2.490000  1.355000 2.775000 2.005000 ;
      RECT 2.735000  0.705000 3.115000 1.035000 ;
      RECT 2.860000  0.365000 3.520000 0.535000 ;
      RECT 2.920000  2.255000 3.670000 2.425000 ;
      RECT 2.945000  1.035000 3.115000 1.415000 ;
      RECT 2.945000  1.415000 3.285000 1.995000 ;
      RECT 3.350000  0.535000 3.520000 0.995000 ;
      RECT 3.350000  0.995000 4.220000 1.165000 ;
      RECT 3.500000  1.165000 4.220000 1.325000 ;
      RECT 3.500000  1.325000 3.670000 2.255000 ;
      RECT 3.760000  0.085000 4.090000 0.825000 ;
      RECT 3.840000  2.135000 4.140000 2.635000 ;
      RECT 3.860000  1.535000 4.580000 1.865000 ;
      RECT 4.360000  0.415000 4.580000 0.825000 ;
      RECT 4.360000  1.865000 4.580000 2.435000 ;
      RECT 4.410000  0.825000 4.580000 0.995000 ;
      RECT 4.410000  0.995000 5.160000 1.325000 ;
      RECT 4.410000  1.325000 4.580000 1.535000 ;
      RECT 4.760000  0.085000 5.045000 0.825000 ;
      RECT 4.760000  1.495000 5.045000 2.635000 ;
      RECT 5.635000  0.085000 5.895000 0.550000 ;
      RECT 5.635000  1.755000 5.895000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.490000  1.785000 2.660000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.950000  1.445000 3.120000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.180000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.720000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.430000 1.755000 2.720000 1.800000 ;
      RECT 2.430000 1.940000 2.720000 1.985000 ;
      RECT 2.890000 1.415000 3.180000 1.460000 ;
      RECT 2.890000 1.600000 3.180000 1.645000 ;
  END
END sky130_fd_sc_hd__dlxtn_2
MACRO sky130_fd_sc_hd__dlxtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.240000 0.415000 5.525000 0.745000 ;
        RECT 5.240000 1.495000 5.525000 2.455000 ;
        RECT 5.355000 0.745000 5.525000 0.995000 ;
        RECT 5.355000 0.995000 6.815000 1.325000 ;
        RECT 5.355000 1.325000 5.525000 1.495000 ;
        RECT 6.115000 0.385000 6.385000 0.995000 ;
        RECT 6.115000 1.325000 6.385000 2.455000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.780000 0.805000 ;
      RECT 0.175000  1.795000 0.780000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 2.005000 ;
      RECT 2.715000  0.705000 3.095000 1.035000 ;
      RECT 2.840000  0.365000 3.500000 0.535000 ;
      RECT 2.900000  2.255000 3.650000 2.425000 ;
      RECT 2.925000  1.035000 3.095000 1.415000 ;
      RECT 2.925000  1.415000 3.265000 1.995000 ;
      RECT 3.330000  0.535000 3.500000 0.995000 ;
      RECT 3.330000  0.995000 4.200000 1.165000 ;
      RECT 3.480000  1.165000 4.200000 1.325000 ;
      RECT 3.480000  1.325000 3.650000 2.255000 ;
      RECT 3.740000  0.085000 4.070000 0.530000 ;
      RECT 3.820000  2.135000 4.120000 2.635000 ;
      RECT 3.840000  1.535000 4.605000 1.865000 ;
      RECT 4.385000  0.415000 4.605000 0.745000 ;
      RECT 4.385000  1.865000 4.605000 2.435000 ;
      RECT 4.435000  0.745000 4.605000 0.995000 ;
      RECT 4.435000  0.995000 5.185000 1.325000 ;
      RECT 4.435000  1.325000 4.605000 1.535000 ;
      RECT 4.785000  0.085000 5.070000 0.715000 ;
      RECT 4.785000  1.495000 5.070000 2.635000 ;
      RECT 5.695000  0.085000 5.945000 0.825000 ;
      RECT 5.695000  1.495000 5.945000 2.635000 ;
      RECT 6.555000  0.085000 6.815000 0.715000 ;
      RECT 6.555000  1.495000 6.815000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.785000 2.640000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.445000 3.100000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 3.160000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 2.700000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.755000 2.700000 1.800000 ;
      RECT 2.410000 1.940000 2.700000 1.985000 ;
      RECT 2.870000 1.415000 3.160000 1.460000 ;
      RECT 2.870000 1.600000 3.160000 1.645000 ;
  END
END sky130_fd_sc_hd__dlxtn_4
MACRO sky130_fd_sc_hd__a221o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855000 1.075000 3.190000 1.105000 ;
        RECT 2.855000 1.105000 4.060000 1.285000 ;
        RECT 3.710000 1.075000 4.060000 1.105000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265000 1.075000 2.680000 1.285000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235000 1.075000 6.035000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.270000 1.075000 7.280000 1.285000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.230000 1.075000 4.725000 1.285000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.735000 1.685000 0.905000 ;
        RECT 0.095000 0.905000 0.325000 1.455000 ;
        RECT 0.095000 1.455000 1.645000 1.625000 ;
        RECT 0.515000 0.255000 0.845000 0.725000 ;
        RECT 0.515000 0.725000 1.685000 0.735000 ;
        RECT 0.555000 1.625000 0.805000 2.465000 ;
        RECT 1.355000 0.255000 1.685000 0.725000 ;
        RECT 1.395000 1.625000 1.645000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.155000  1.795000 0.385000 2.635000 ;
      RECT 0.175000  0.085000 0.345000 0.555000 ;
      RECT 0.495000  1.075000 1.845000 1.115000 ;
      RECT 0.495000  1.115000 1.985000 1.285000 ;
      RECT 0.975000  1.795000 1.225000 2.635000 ;
      RECT 1.015000  0.085000 1.185000 0.555000 ;
      RECT 1.815000  1.285000 1.985000 1.455000 ;
      RECT 1.815000  1.455000 5.065000 1.625000 ;
      RECT 1.815000  1.795000 2.065000 2.635000 ;
      RECT 1.855000  0.085000 2.025000 0.555000 ;
      RECT 1.855000  0.735000 2.525000 0.905000 ;
      RECT 1.945000  0.905000 2.165000 0.935000 ;
      RECT 2.195000  0.255000 2.525000 0.735000 ;
      RECT 2.235000  1.795000 4.230000 1.875000 ;
      RECT 2.235000  1.875000 5.575000 1.965000 ;
      RECT 2.235000  1.965000 2.485000 2.465000 ;
      RECT 2.655000  2.135000 2.905000 2.635000 ;
      RECT 2.695000  0.085000 2.865000 0.895000 ;
      RECT 3.075000  1.965000 3.330000 2.465000 ;
      RECT 3.080000  0.305000 4.305000 0.475000 ;
      RECT 3.190000  0.735000 3.885000 0.905000 ;
      RECT 3.315000  0.905000 3.610000 0.935000 ;
      RECT 3.500000  2.135000 3.750000 2.635000 ;
      RECT 3.550000  0.645000 3.885000 0.735000 ;
      RECT 3.940000  2.215000 6.385000 2.295000 ;
      RECT 3.940000  2.295000 7.225000 2.465000 ;
      RECT 4.055000  0.475000 4.305000 0.725000 ;
      RECT 4.055000  0.725000 5.065000 0.905000 ;
      RECT 4.060000  1.965000 5.575000 2.045000 ;
      RECT 4.405000  1.625000 4.735000 1.705000 ;
      RECT 4.475000  0.085000 4.645000 0.555000 ;
      RECT 4.815000  0.255000 5.985000 0.475000 ;
      RECT 4.815000  0.475000 5.065000 0.725000 ;
      RECT 4.895000  0.905000 5.065000 1.455000 ;
      RECT 5.235000  0.645000 6.505000 0.725000 ;
      RECT 5.235000  0.725000 7.345000 0.905000 ;
      RECT 5.245000  1.455000 6.805000 1.625000 ;
      RECT 5.245000  1.625000 5.575000 1.875000 ;
      RECT 5.745000  1.795000 6.385000 2.215000 ;
      RECT 6.555000  1.625000 6.805000 2.125000 ;
      RECT 6.675000  0.085000 6.845000 0.555000 ;
      RECT 6.975000  1.785000 7.225000 2.295000 ;
      RECT 7.015000  0.255000 7.345000 0.725000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 1.995000  0.765000 2.165000 0.935000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.400000  0.765000 3.570000 0.935000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 1.935000 0.735000 2.225000 0.780000 ;
      RECT 1.935000 0.780000 3.630000 0.920000 ;
      RECT 1.935000 0.920000 2.225000 0.965000 ;
      RECT 3.340000 0.735000 3.630000 0.780000 ;
      RECT 3.340000 0.920000 3.630000 0.965000 ;
  END
END sky130_fd_sc_hd__a221o_4
MACRO sky130_fd_sc_hd__a221o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 0.675000 2.255000 1.075000 ;
        RECT 1.970000 1.075000 2.300000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 1.075000 2.835000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 1.075000 1.700000 1.275000 ;
        RECT 1.420000 0.675000 1.700000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.075000 1.055000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.440000 1.285000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.320000 0.255000 3.575000 0.585000 ;
        RECT 3.320000 1.795000 3.575000 2.465000 ;
        RECT 3.390000 0.585000 3.575000 0.665000 ;
        RECT 3.405000 0.665000 3.575000 1.795000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.735000 ;
      RECT 0.175000  0.735000 1.240000 0.905000 ;
      RECT 0.175000  1.455000 3.235000 1.625000 ;
      RECT 0.175000  1.625000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.565000 ;
      RECT 0.515000  1.795000 0.845000 2.295000 ;
      RECT 0.515000  2.295000 1.685000 2.465000 ;
      RECT 1.015000  1.795000 2.650000 2.035000 ;
      RECT 1.015000  2.035000 1.245000 2.125000 ;
      RECT 1.070000  0.255000 2.605000 0.505000 ;
      RECT 1.070000  0.505000 1.240000 0.735000 ;
      RECT 1.355000  2.255000 1.685000 2.295000 ;
      RECT 1.875000  2.215000 2.230000 2.635000 ;
      RECT 2.400000  2.035000 2.650000 2.465000 ;
      RECT 2.435000  0.505000 2.605000 0.735000 ;
      RECT 2.435000  0.735000 3.235000 0.905000 ;
      RECT 2.775000  0.085000 3.105000 0.565000 ;
      RECT 2.820000  1.875000 3.150000 2.635000 ;
      RECT 3.065000  0.905000 3.235000 1.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a221o_1
MACRO sky130_fd_sc_hd__a221o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 0.675000 2.255000 1.075000 ;
        RECT 1.970000 1.075000 2.300000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 1.075000 2.835000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 1.075000 1.700000 1.275000 ;
        RECT 1.420000 0.675000 1.700000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.075000 1.055000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.440000 1.285000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.320000 0.255000 3.575000 0.585000 ;
        RECT 3.320000 1.795000 3.575000 2.465000 ;
        RECT 3.390000 0.585000 3.575000 0.665000 ;
        RECT 3.405000 0.665000 3.575000 1.795000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.735000 ;
      RECT 0.175000  0.735000 1.240000 0.905000 ;
      RECT 0.175000  1.455000 3.235000 1.625000 ;
      RECT 0.175000  1.625000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.565000 ;
      RECT 0.515000  1.795000 0.845000 2.295000 ;
      RECT 0.515000  2.295000 1.685000 2.465000 ;
      RECT 1.015000  1.795000 2.650000 2.035000 ;
      RECT 1.015000  2.035000 1.245000 2.125000 ;
      RECT 1.070000  0.255000 2.605000 0.505000 ;
      RECT 1.070000  0.505000 1.240000 0.735000 ;
      RECT 1.355000  2.255000 1.685000 2.295000 ;
      RECT 1.875000  2.215000 2.230000 2.635000 ;
      RECT 2.400000  2.035000 2.650000 2.465000 ;
      RECT 2.435000  0.505000 2.605000 0.735000 ;
      RECT 2.435000  0.735000 3.235000 0.905000 ;
      RECT 2.775000  0.085000 3.105000 0.565000 ;
      RECT 2.820000  1.875000 3.150000 2.635000 ;
      RECT 3.065000  0.905000 3.235000 1.455000 ;
      RECT 3.745000  0.085000 3.915000 0.980000 ;
      RECT 3.745000  1.445000 3.915000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a221o_2
MACRO sky130_fd_sc_hd__or2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 2.085000 1.730000 2.415000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.325000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.400000 0.415000 2.630000 0.760000 ;
        RECT 2.400000 1.495000 2.630000 2.465000 ;
        RECT 2.460000 0.760000 2.630000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.105000  0.265000 0.420000 0.735000 ;
      RECT 0.105000  0.735000 0.840000 0.905000 ;
      RECT 0.590000  0.085000 1.320000 0.565000 ;
      RECT 0.595000  0.905000 0.840000 0.995000 ;
      RECT 0.595000  0.995000 1.330000 1.325000 ;
      RECT 0.595000  1.325000 0.765000 1.885000 ;
      RECT 0.985000  1.495000 2.230000 1.665000 ;
      RECT 0.985000  1.665000 1.405000 1.915000 ;
      RECT 1.490000  0.305000 1.660000 0.655000 ;
      RECT 1.490000  0.655000 2.230000 0.825000 ;
      RECT 1.830000  0.085000 2.210000 0.485000 ;
      RECT 1.910000  1.835000 2.190000 2.635000 ;
      RECT 2.060000  0.825000 2.230000 0.995000 ;
      RECT 2.060000  0.995000 2.290000 1.325000 ;
      RECT 2.060000  1.325000 2.230000 1.495000 ;
      RECT 2.800000  0.085000 3.055000 0.925000 ;
      RECT 2.800000  1.460000 3.055000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__or2b_2
MACRO sky130_fd_sc_hd__or2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.630000 1.075000 2.320000 1.275000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.955000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 0.290000 2.655000 0.735000 ;
        RECT 2.325000 0.735000 4.055000 0.905000 ;
        RECT 2.365000 1.785000 3.455000 1.955000 ;
        RECT 2.365000 1.955000 2.615000 2.465000 ;
        RECT 2.830000 1.445000 4.055000 1.615000 ;
        RECT 2.830000 1.615000 3.455000 1.785000 ;
        RECT 3.165000 0.290000 3.495000 0.735000 ;
        RECT 3.205000 1.955000 3.455000 2.465000 ;
        RECT 3.670000 0.905000 4.055000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  2.125000 0.345000 2.635000 ;
      RECT 0.110000  0.265000 0.420000 0.735000 ;
      RECT 0.110000  0.735000 0.845000 0.905000 ;
      RECT 0.590000  0.085000 1.245000 0.565000 ;
      RECT 0.595000  0.905000 0.845000 0.995000 ;
      RECT 0.595000  0.995000 1.120000 1.325000 ;
      RECT 0.595000  1.325000 0.765000 2.465000 ;
      RECT 0.990000  1.495000 2.660000 1.615000 ;
      RECT 0.990000  1.615000 1.460000 2.465000 ;
      RECT 1.290000  0.735000 1.745000 0.905000 ;
      RECT 1.290000  0.905000 1.460000 1.445000 ;
      RECT 1.290000  1.445000 2.660000 1.495000 ;
      RECT 1.415000  0.305000 1.745000 0.735000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
      RECT 1.980000  0.085000 2.155000 0.905000 ;
      RECT 2.490000  1.075000 3.500000 1.245000 ;
      RECT 2.490000  1.245000 2.660000 1.445000 ;
      RECT 2.785000  2.135000 3.035000 2.635000 ;
      RECT 2.825000  0.085000 2.995000 0.550000 ;
      RECT 3.625000  1.795000 3.875000 2.635000 ;
      RECT 3.665000  0.085000 3.835000 0.550000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__or2b_4
MACRO sky130_fd_sc_hd__or2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 2.085000 1.735000 2.415000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.325000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 0.415000 2.675000 0.760000 ;
        RECT 2.405000 1.495000 2.675000 2.465000 ;
        RECT 2.505000 0.760000 2.675000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.110000  0.265000 0.420000 0.735000 ;
      RECT 0.110000  0.735000 0.845000 0.905000 ;
      RECT 0.590000  0.085000 1.325000 0.565000 ;
      RECT 0.595000  0.905000 0.845000 0.995000 ;
      RECT 0.595000  0.995000 1.335000 1.325000 ;
      RECT 0.595000  1.325000 0.765000 1.885000 ;
      RECT 0.990000  1.495000 2.235000 1.665000 ;
      RECT 0.990000  1.665000 1.410000 1.915000 ;
      RECT 1.495000  0.305000 1.665000 0.655000 ;
      RECT 1.495000  0.655000 2.235000 0.825000 ;
      RECT 1.835000  0.085000 2.215000 0.485000 ;
      RECT 1.915000  1.835000 2.195000 2.635000 ;
      RECT 2.065000  0.825000 2.235000 0.995000 ;
      RECT 2.065000  0.995000 2.295000 1.325000 ;
      RECT 2.065000  1.325000 2.235000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__or2b_1
MACRO sky130_fd_sc_hd__o211a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.300000 1.075000 1.720000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.890000 1.075000 2.220000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.390000 1.075000 2.720000 1.275000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.245000 1.075000 3.595000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.425000 0.885000 ;
        RECT 0.085000 0.885000 0.260000 1.495000 ;
        RECT 0.085000 1.495000 0.425000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.430000  1.075000 1.125000 1.245000 ;
      RECT 0.595000  0.085000 0.845000 0.885000 ;
      RECT 0.595000  1.495000 0.765000 2.635000 ;
      RECT 0.955000  1.245000 1.125000 1.495000 ;
      RECT 0.955000  1.495000 3.390000 1.665000 ;
      RECT 1.035000  0.255000 1.365000 0.735000 ;
      RECT 1.035000  0.735000 2.260000 0.905000 ;
      RECT 1.035000  1.835000 1.285000 2.635000 ;
      RECT 1.535000  0.085000 1.760000 0.545000 ;
      RECT 1.930000  0.255000 2.260000 0.735000 ;
      RECT 1.930000  1.665000 2.260000 2.465000 ;
      RECT 2.560000  1.835000 2.890000 2.635000 ;
      RECT 2.890000  0.255000 3.390000 0.865000 ;
      RECT 2.890000  0.865000 3.060000 1.495000 ;
      RECT 3.060000  1.665000 3.390000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o211a_1
MACRO sky130_fd_sc_hd__o211a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.490000 1.035000 4.845000 1.495000 ;
        RECT 4.490000 1.495000 6.290000 1.685000 ;
        RECT 5.890000 1.035000 6.290000 1.495000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.030000 1.035000 5.705000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.540000 0.995000 2.830000 1.445000 ;
        RECT 2.540000 1.445000 4.280000 1.685000 ;
        RECT 3.950000 1.035000 4.280000 1.445000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.055000 1.035000 3.740000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.911000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.635000 1.605000 0.805000 ;
        RECT 0.085000 0.805000 0.365000 1.435000 ;
        RECT 0.085000 1.435000 2.030000 1.700000 ;
        RECT 0.595000 0.255000 0.765000 0.615000 ;
        RECT 0.595000 0.615000 1.605000 0.635000 ;
        RECT 0.980000 1.700000 1.160000 2.465000 ;
        RECT 1.435000 0.255000 1.605000 0.615000 ;
        RECT 1.840000 1.700000 2.030000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.480000  1.870000 0.810000 2.635000 ;
      RECT 0.535000  1.065000 2.370000 1.265000 ;
      RECT 0.935000  0.085000 1.265000 0.445000 ;
      RECT 1.340000  1.870000 1.670000 2.635000 ;
      RECT 1.775000  0.085000 2.140000 0.465000 ;
      RECT 2.200000  0.635000 3.520000 0.815000 ;
      RECT 2.200000  0.815000 2.370000 1.065000 ;
      RECT 2.200000  1.265000 2.370000 1.855000 ;
      RECT 2.200000  1.855000 5.485000 2.025000 ;
      RECT 2.200000  2.200000 2.530000 2.635000 ;
      RECT 2.330000  0.255000 4.500000 0.465000 ;
      RECT 2.700000  2.025000 3.060000 2.465000 ;
      RECT 3.285000  2.195000 3.615000 2.635000 ;
      RECT 3.785000  2.025000 4.120000 2.465000 ;
      RECT 4.170000  0.465000 4.500000 0.695000 ;
      RECT 4.170000  0.695000 6.345000 0.865000 ;
      RECT 4.290000  2.195000 4.555000 2.635000 ;
      RECT 4.670000  0.085000 4.985000 0.525000 ;
      RECT 5.155000  0.255000 5.485000 0.695000 ;
      RECT 5.155000  2.025000 5.485000 2.465000 ;
      RECT 5.655000  0.085000 5.845000 0.525000 ;
      RECT 6.015000  0.255000 6.345000 0.695000 ;
      RECT 6.015000  1.915000 6.345000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__o211a_4
MACRO sky130_fd_sc_hd__o211a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 0.995000 2.325000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.995000 1.820000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.880000 0.995000 1.240000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.360000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.720000 0.255000 3.050000 0.615000 ;
        RECT 2.720000 0.615000 3.540000 0.785000 ;
        RECT 2.810000 1.905000 3.540000 2.075000 ;
        RECT 2.810000 2.075000 3.000000 2.465000 ;
        RECT 3.345000 0.785000 3.540000 1.905000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  1.510000 2.665000 1.765000 ;
      RECT 0.090000  1.765000 0.355000 2.465000 ;
      RECT 0.095000  0.255000 0.430000 0.425000 ;
      RECT 0.095000  0.425000 0.710000 0.825000 ;
      RECT 0.525000  1.935000 0.855000 2.635000 ;
      RECT 0.530000  0.825000 0.710000 1.510000 ;
      RECT 0.880000  0.635000 2.150000 0.825000 ;
      RECT 1.025000  1.765000 1.695000 2.465000 ;
      RECT 1.390000  0.085000 1.725000 0.465000 ;
      RECT 2.200000  1.935000 2.630000 2.635000 ;
      RECT 2.315000  0.085000 2.550000 0.525000 ;
      RECT 2.495000  0.995000 3.175000 1.325000 ;
      RECT 2.495000  1.325000 2.665000 1.510000 ;
      RECT 3.170000  2.255000 3.500000 2.635000 ;
      RECT 3.220000  0.085000 3.550000 0.445000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o211a_2
MACRO sky130_fd_sc_hd__nor4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 1.075000 1.805000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.075000 3.750000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.985000 1.075000 5.685000 1.285000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.810000 1.075000 8.655000 1.285000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.845000 0.725000 ;
        RECT 0.515000 0.725000 7.245000 0.905000 ;
        RECT 1.355000 0.255000 1.685000 0.725000 ;
        RECT 2.195000 0.255000 2.525000 0.725000 ;
        RECT 3.035000 0.255000 3.365000 0.725000 ;
        RECT 4.395000 0.255000 4.725000 0.725000 ;
        RECT 5.235000 0.255000 5.565000 0.725000 ;
        RECT 6.075000 0.255000 6.405000 0.725000 ;
        RECT 6.115000 0.905000 6.465000 1.455000 ;
        RECT 6.115000 1.455000 7.205000 1.625000 ;
        RECT 6.115000 1.625000 6.365000 2.125000 ;
        RECT 6.915000 0.255000 7.245000 0.725000 ;
        RECT 6.955000 1.625000 7.205000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.095000  1.455000 2.065000 1.625000 ;
      RECT 0.095000  1.625000 0.425000 2.465000 ;
      RECT 0.175000  0.085000 0.345000 0.895000 ;
      RECT 0.595000  1.795000 0.805000 2.635000 ;
      RECT 0.975000  1.625000 1.225000 2.465000 ;
      RECT 1.015000  0.085000 1.185000 0.555000 ;
      RECT 1.395000  1.795000 1.645000 2.635000 ;
      RECT 1.815000  1.625000 2.065000 2.295000 ;
      RECT 1.815000  2.295000 3.745000 2.465000 ;
      RECT 1.855000  0.085000 2.025000 0.555000 ;
      RECT 2.235000  1.455000 5.525000 1.625000 ;
      RECT 2.235000  1.625000 2.485000 2.125000 ;
      RECT 2.655000  1.795000 2.905000 2.295000 ;
      RECT 2.695000  0.085000 2.865000 0.555000 ;
      RECT 3.075000  1.625000 3.325000 2.125000 ;
      RECT 3.495000  1.795000 3.745000 2.295000 ;
      RECT 3.535000  0.085000 4.225000 0.555000 ;
      RECT 4.015000  1.795000 4.265000 2.295000 ;
      RECT 4.015000  2.295000 7.625000 2.465000 ;
      RECT 4.435000  1.625000 4.685000 2.125000 ;
      RECT 4.855000  1.795000 5.105000 2.295000 ;
      RECT 4.895000  0.085000 5.065000 0.555000 ;
      RECT 5.275000  1.625000 5.525000 2.125000 ;
      RECT 5.695000  1.455000 5.945000 2.295000 ;
      RECT 5.735000  0.085000 5.905000 0.555000 ;
      RECT 6.535000  1.795000 6.785000 2.295000 ;
      RECT 6.575000  0.085000 6.745000 0.555000 ;
      RECT 6.635000  1.075000 7.640000 1.285000 ;
      RECT 7.375000  1.795000 7.625000 2.295000 ;
      RECT 7.415000  0.085000 7.585000 0.555000 ;
      RECT 7.470000  0.735000 8.185000 0.905000 ;
      RECT 7.470000  0.905000 7.640000 1.075000 ;
      RECT 7.470000  1.285000 7.640000 1.455000 ;
      RECT 7.470000  1.455000 8.185000 1.625000 ;
      RECT 7.810000  0.255000 8.185000 0.735000 ;
      RECT 7.850000  1.625000 8.185000 2.465000 ;
      RECT 8.355000  0.085000 8.585000 0.905000 ;
      RECT 8.355000  1.455000 8.585000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4b_4
MACRO sky130_fd_sc_hd__nor4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 0.995000 2.275000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.995000 1.785000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 0.995000 1.285000 1.615000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.995000 2.795000 1.615000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.871000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.655000 1.925000 0.825000 ;
        RECT 0.085000 0.825000 0.345000 2.450000 ;
        RECT 0.855000 0.300000 1.055000 0.655000 ;
        RECT 1.725000 0.310000 1.925000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.355000  0.085000 0.685000 0.480000 ;
      RECT 0.525000  0.995000 0.745000 1.795000 ;
      RECT 0.525000  1.795000 3.135000 2.005000 ;
      RECT 1.225000  0.085000 1.555000 0.485000 ;
      RECT 2.095000  0.085000 2.425000 0.825000 ;
      RECT 2.095000  2.185000 2.425000 2.635000 ;
      RECT 2.660000  0.405000 2.830000 0.655000 ;
      RECT 2.660000  0.655000 3.135000 0.825000 ;
      RECT 2.965000  0.825000 3.135000 1.795000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4b_1
MACRO sky130_fd_sc_hd__nor4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 1.240000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 1.075000 2.635000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815000 1.075000 3.535000 1.285000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.805000 1.075000 5.435000 1.285000 ;
        RECT 5.185000 1.285000 5.435000 1.955000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.255000 0.845000 0.725000 ;
        RECT 0.515000 0.725000 3.920000 0.905000 ;
        RECT 1.355000 0.255000 1.685000 0.725000 ;
        RECT 2.750000 0.255000 3.080000 0.725000 ;
        RECT 3.590000 0.255000 3.920000 0.725000 ;
        RECT 3.630000 1.455000 4.035000 1.625000 ;
        RECT 3.630000 1.625000 3.880000 2.125000 ;
        RECT 3.715000 0.905000 3.920000 1.075000 ;
        RECT 3.715000 1.075000 4.035000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.905000 ;
      RECT 0.085000  1.455000 2.105000 1.625000 ;
      RECT 0.085000  1.625000 0.425000 2.465000 ;
      RECT 0.595000  1.795000 0.805000 2.635000 ;
      RECT 0.975000  1.625000 1.225000 2.465000 ;
      RECT 1.015000  0.085000 1.185000 0.555000 ;
      RECT 1.395000  1.795000 1.605000 2.295000 ;
      RECT 1.395000  2.295000 3.040000 2.465000 ;
      RECT 1.775000  1.625000 2.105000 2.125000 ;
      RECT 1.855000  0.085000 2.580000 0.555000 ;
      RECT 2.275000  1.455000 3.460000 1.625000 ;
      RECT 2.275000  1.625000 2.660000 2.125000 ;
      RECT 2.830000  1.795000 3.040000 2.295000 ;
      RECT 3.210000  1.625000 3.460000 2.295000 ;
      RECT 3.210000  2.295000 4.295000 2.465000 ;
      RECT 3.250000  0.085000 3.420000 0.555000 ;
      RECT 4.050000  1.795000 4.295000 2.295000 ;
      RECT 4.090000  0.085000 4.295000 0.895000 ;
      RECT 4.320000  1.075000 4.635000 1.245000 ;
      RECT 4.465000  0.380000 4.820000 0.905000 ;
      RECT 4.465000  0.905000 4.635000 1.075000 ;
      RECT 4.465000  1.245000 4.635000 2.035000 ;
      RECT 4.465000  2.035000 4.820000 2.450000 ;
      RECT 4.990000  0.085000 5.240000 0.825000 ;
      RECT 4.990000  2.135000 5.240000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4b_2
MACRO sky130_fd_sc_hd__ebufn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 0.765000 0.780000 1.675000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.811500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.765000 1.280000 1.425000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 1.445000 5.895000 1.725000 ;
        RECT 4.145000 0.615000 5.895000 0.855000 ;
        RECT 5.675000 0.855000 5.895000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.280000 0.345000 0.665000 ;
      RECT 0.085000  0.665000 0.320000 1.765000 ;
      RECT 0.085000  1.765000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.930000 0.595000 ;
      RECT 0.515000  1.845000 0.930000 2.635000 ;
      RECT 1.100000  0.255000 1.725000 0.595000 ;
      RECT 1.100000  1.595000 1.725000 1.765000 ;
      RECT 1.100000  1.765000 1.355000 2.465000 ;
      RECT 1.450000  0.595000 1.725000 1.025000 ;
      RECT 1.450000  1.025000 3.810000 1.275000 ;
      RECT 1.450000  1.275000 1.725000 1.595000 ;
      RECT 1.565000  1.935000 5.895000 2.105000 ;
      RECT 1.565000  2.105000 1.810000 2.465000 ;
      RECT 1.895000  0.255000 2.175000 0.655000 ;
      RECT 1.895000  0.655000 3.975000 0.855000 ;
      RECT 1.895000  1.895000 5.895000 1.935000 ;
      RECT 1.980000  2.275000 2.310000 2.635000 ;
      RECT 2.345000  0.085000 2.675000 0.485000 ;
      RECT 2.480000  2.105000 2.650000 2.465000 ;
      RECT 2.820000  2.275000 3.150000 2.635000 ;
      RECT 2.845000  0.275000 3.015000 0.655000 ;
      RECT 3.185000  0.085000 3.515000 0.485000 ;
      RECT 3.320000  2.105000 5.895000 2.465000 ;
      RECT 3.685000  0.255000 5.735000 0.445000 ;
      RECT 3.685000  0.445000 3.975000 0.655000 ;
      RECT 3.980000  1.025000 5.505000 1.275000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.150000  1.105000 0.320000 1.275000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.310000  1.105000 4.480000 1.275000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 0.085000 1.075000 0.380000 1.120000 ;
      RECT 0.085000 1.120000 4.540000 1.260000 ;
      RECT 0.085000 1.260000 0.380000 1.305000 ;
      RECT 4.250000 1.075000 4.540000 1.120000 ;
      RECT 4.250000 1.260000 4.540000 1.305000 ;
  END
END sky130_fd_sc_hd__ebufn_4
MACRO sky130_fd_sc_hd__ebufn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.355000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.309000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 1.075000 1.240000 1.630000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.601000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.495000 3.595000 2.465000 ;
        RECT 3.125000 0.255000 3.595000 0.825000 ;
        RECT 3.255000 0.825000 3.595000 1.495000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.280000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.185000 0.825000 ;
      RECT 0.085000  1.785000 0.740000 2.005000 ;
      RECT 0.085000  2.005000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.445000 ;
      RECT 0.515000  2.175000 0.845000 2.635000 ;
      RECT 0.525000  0.825000 0.740000 1.785000 ;
      RECT 1.015000  0.255000 2.025000 0.465000 ;
      RECT 1.015000  0.465000 1.185000 0.615000 ;
      RECT 1.015000  1.800000 1.805000 2.005000 ;
      RECT 1.015000  2.005000 1.270000 2.460000 ;
      RECT 1.355000  0.635000 1.685000 0.885000 ;
      RECT 1.410000  0.885000 1.685000 1.075000 ;
      RECT 1.410000  1.075000 2.535000 1.325000 ;
      RECT 1.410000  1.325000 1.805000 1.800000 ;
      RECT 1.440000  2.175000 1.805000 2.635000 ;
      RECT 1.855000  0.465000 2.025000 0.735000 ;
      RECT 1.855000  0.735000 2.955000 0.905000 ;
      RECT 2.195000  0.085000 2.955000 0.565000 ;
      RECT 2.705000  0.905000 2.955000 0.995000 ;
      RECT 2.705000  0.995000 3.085000 1.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__ebufn_1
MACRO sky130_fd_sc_hd__ebufn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 0.765000 0.780000 1.675000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.441000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.765000 1.280000 1.275000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.905000 1.445000 4.055000 1.625000 ;
        RECT 1.905000 1.625000 3.625000 1.765000 ;
        RECT 3.295000 0.635000 4.055000 0.855000 ;
        RECT 3.295000 1.765000 3.625000 2.125000 ;
        RECT 3.825000 0.855000 4.055000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.280000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 0.320000 1.845000 ;
      RECT 0.085000  1.845000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.850000 0.595000 ;
      RECT 0.515000  1.845000 0.950000 2.635000 ;
      RECT 1.020000  0.255000 1.730000 0.595000 ;
      RECT 1.120000  1.445000 1.735000 1.765000 ;
      RECT 1.120000  1.765000 1.410000 2.465000 ;
      RECT 1.450000  0.595000 1.730000 1.025000 ;
      RECT 1.450000  1.025000 2.965000 1.275000 ;
      RECT 1.450000  1.275000 1.735000 1.445000 ;
      RECT 1.600000  1.935000 3.125000 2.105000 ;
      RECT 1.600000  2.105000 1.810000 2.465000 ;
      RECT 1.900000  0.255000 2.170000 0.655000 ;
      RECT 1.900000  0.655000 3.125000 0.855000 ;
      RECT 1.980000  2.275000 2.310000 2.635000 ;
      RECT 2.340000  0.085000 2.670000 0.485000 ;
      RECT 2.480000  2.105000 3.125000 2.295000 ;
      RECT 2.480000  2.295000 4.055000 2.465000 ;
      RECT 2.840000  0.275000 4.050000 0.465000 ;
      RECT 2.840000  0.465000 3.125000 0.655000 ;
      RECT 3.245000  1.025000 3.655000 1.275000 ;
      RECT 3.795000  1.795000 4.055000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.150000  1.105000 0.320000 1.275000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.380000  1.105000 3.550000 1.275000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
    LAYER met1 ;
      RECT 0.085000 1.075000 0.380000 1.120000 ;
      RECT 0.085000 1.120000 3.610000 1.260000 ;
      RECT 0.085000 1.260000 0.380000 1.305000 ;
      RECT 3.320000 1.075000 3.610000 1.120000 ;
      RECT 3.320000 1.260000 3.610000 1.305000 ;
  END
END sky130_fd_sc_hd__ebufn_2
MACRO sky130_fd_sc_hd__ebufn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.430000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.375500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.970000 0.620000 1.305000 0.995000 ;
        RECT 0.970000 0.995000 1.430000 1.325000 ;
        RECT 0.970000 1.325000 1.305000 1.695000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.445000 9.575000 1.725000 ;
        RECT 6.275000 0.615000 9.575000 0.855000 ;
        RECT 9.325000 0.855000 9.575000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.085000  0.085000 0.445000 0.825000 ;
      RECT 0.085000  1.785000 0.445000 2.635000 ;
      RECT 0.600000  0.995000 0.800000 1.615000 ;
      RECT 0.615000  0.280000 0.800000 0.995000 ;
      RECT 0.615000  1.615000 0.800000 2.465000 ;
      RECT 0.970000  0.085000 1.305000 0.445000 ;
      RECT 0.970000  1.865000 1.305000 2.635000 ;
      RECT 1.475000  0.255000 1.985000 0.825000 ;
      RECT 1.475000  1.495000 1.825000 2.465000 ;
      RECT 1.600000  0.825000 1.985000 1.025000 ;
      RECT 1.600000  1.025000 5.925000 1.275000 ;
      RECT 1.600000  1.275000 1.825000 1.495000 ;
      RECT 1.995000  1.895000 9.575000 2.065000 ;
      RECT 1.995000  2.065000 2.245000 2.465000 ;
      RECT 2.155000  0.255000 2.485000 0.655000 ;
      RECT 2.155000  0.655000 6.105000 0.855000 ;
      RECT 2.415000  2.235000 2.745000 2.635000 ;
      RECT 2.655000  0.085000 2.985000 0.485000 ;
      RECT 2.915000  2.065000 3.085000 2.465000 ;
      RECT 3.155000  0.275000 3.325000 0.655000 ;
      RECT 3.255000  2.235000 3.585000 2.635000 ;
      RECT 3.495000  0.085000 3.825000 0.485000 ;
      RECT 3.755000  2.065000 3.925000 2.465000 ;
      RECT 3.995000  0.255000 4.165000 0.655000 ;
      RECT 4.095000  2.235000 4.425000 2.635000 ;
      RECT 4.335000  0.085000 4.665000 0.485000 ;
      RECT 4.595000  2.065000 4.765000 2.465000 ;
      RECT 4.835000  0.275000 5.005000 0.655000 ;
      RECT 4.935000  2.235000 5.265000 2.635000 ;
      RECT 5.175000  0.085000 5.505000 0.485000 ;
      RECT 5.435000  2.065000 9.575000 2.465000 ;
      RECT 5.675000  0.255000 9.575000 0.445000 ;
      RECT 5.675000  0.445000 6.105000 0.655000 ;
      RECT 6.175000  1.025000 9.155000 1.275000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  1.105000 0.775000 1.275000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.580000  1.105000 6.750000 1.275000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.545000 1.075000 0.835000 1.120000 ;
      RECT 0.545000 1.120000 6.810000 1.260000 ;
      RECT 0.545000 1.260000 0.835000 1.305000 ;
      RECT 6.520000 1.075000 6.810000 1.120000 ;
      RECT 6.520000 1.260000 6.810000 1.305000 ;
  END
END sky130_fd_sc_hd__ebufn_8
MACRO sky130_fd_sc_hd__dfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.370000 0.715000 1.650000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.890000 1.495000 7.300000 1.575000 ;
        RECT 6.890000 1.575000 7.220000 2.420000 ;
        RECT 6.900000 0.305000 7.230000 0.740000 ;
        RECT 6.900000 0.740000 7.300000 0.825000 ;
        RECT 7.055000 0.825000 7.300000 0.865000 ;
        RECT 7.065000 1.445000 7.300000 1.495000 ;
        RECT 7.110000 0.865000 7.300000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.810000 1.495000 9.145000 2.465000 ;
        RECT 8.890000 0.265000 9.145000 0.885000 ;
        RECT 8.930000 0.885000 9.145000 1.495000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.200000 2.465000 ;
      RECT 1.440000  2.175000 1.705000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.820000  0.675000 2.045000 0.805000 ;
      RECT 1.820000  0.805000 1.990000 1.910000 ;
      RECT 1.820000  1.910000 2.125000 2.040000 ;
      RECT 1.875000  0.365000 2.210000 0.535000 ;
      RECT 1.875000  0.535000 2.045000 0.675000 ;
      RECT 1.875000  2.040000 2.125000 2.465000 ;
      RECT 2.160000  1.125000 2.400000 1.720000 ;
      RECT 2.215000  0.735000 2.740000 0.955000 ;
      RECT 2.335000  2.190000 3.440000 2.360000 ;
      RECT 2.405000  0.365000 3.080000 0.535000 ;
      RECT 2.570000  0.955000 2.740000 1.655000 ;
      RECT 2.570000  1.655000 3.100000 2.020000 ;
      RECT 2.910000  0.535000 3.080000 1.315000 ;
      RECT 2.910000  1.315000 3.780000 1.485000 ;
      RECT 3.270000  1.485000 3.780000 1.575000 ;
      RECT 3.270000  1.575000 3.440000 2.190000 ;
      RECT 3.290000  0.765000 4.120000 1.065000 ;
      RECT 3.290000  1.065000 3.490000 1.095000 ;
      RECT 3.400000  0.085000 3.770000 0.585000 ;
      RECT 3.610000  1.245000 3.780000 1.315000 ;
      RECT 3.610000  1.835000 3.780000 2.635000 ;
      RECT 3.950000  0.365000 4.355000 0.535000 ;
      RECT 3.950000  0.535000 4.120000 0.765000 ;
      RECT 3.950000  1.065000 4.120000 2.135000 ;
      RECT 3.950000  2.135000 4.200000 2.465000 ;
      RECT 4.290000  1.245000 4.480000 1.965000 ;
      RECT 4.425000  2.165000 5.310000 2.335000 ;
      RECT 4.505000  0.705000 4.970000 1.035000 ;
      RECT 4.525000  0.365000 5.310000 0.535000 ;
      RECT 4.650000  1.035000 4.970000 1.995000 ;
      RECT 5.140000  0.535000 5.310000 0.995000 ;
      RECT 5.140000  0.995000 6.020000 1.325000 ;
      RECT 5.140000  1.325000 5.310000 2.165000 ;
      RECT 5.480000  1.530000 6.380000 1.905000 ;
      RECT 5.490000  2.135000 5.805000 2.635000 ;
      RECT 5.585000  0.085000 5.795000 0.615000 ;
      RECT 6.040000  1.905000 6.380000 2.465000 ;
      RECT 6.060000  0.300000 6.390000 0.825000 ;
      RECT 6.190000  0.825000 6.390000 0.995000 ;
      RECT 6.190000  0.995000 6.940000 1.325000 ;
      RECT 6.190000  1.325000 6.380000 1.530000 ;
      RECT 6.550000  1.625000 6.720000 2.635000 ;
      RECT 6.560000  0.085000 6.730000 0.695000 ;
      RECT 7.390000  1.720000 7.565000 2.635000 ;
      RECT 7.400000  0.085000 7.570000 0.600000 ;
      RECT 7.905000  0.345000 8.165000 0.615000 ;
      RECT 7.905000  1.715000 8.235000 2.445000 ;
      RECT 7.965000  0.615000 8.165000 0.995000 ;
      RECT 7.965000  0.995000 8.760000 1.325000 ;
      RECT 7.965000  1.325000 8.235000 1.715000 ;
      RECT 8.390000  0.085000 8.720000 0.825000 ;
      RECT 8.425000  1.495000 8.640000 2.635000 ;
      RECT 9.315000  0.085000 9.565000 0.905000 ;
      RECT 9.315000  1.495000 9.565000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.630000  1.785000 0.800000 1.955000 ;
      RECT 1.025000  1.445000 1.195000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.215000  1.445000 2.385000 1.615000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.730000  1.785000 2.900000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.300000  1.785000 4.470000 1.955000 ;
      RECT 4.735000  1.445000 4.905000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.570000 1.755000 0.860000 1.800000 ;
      RECT 0.570000 1.800000 4.530000 1.940000 ;
      RECT 0.570000 1.940000 0.860000 1.985000 ;
      RECT 0.965000 1.415000 1.255000 1.460000 ;
      RECT 0.965000 1.460000 4.965000 1.600000 ;
      RECT 0.965000 1.600000 1.255000 1.645000 ;
      RECT 2.155000 1.415000 2.445000 1.460000 ;
      RECT 2.155000 1.600000 2.445000 1.645000 ;
      RECT 2.670000 1.755000 2.960000 1.800000 ;
      RECT 2.670000 1.940000 2.960000 1.985000 ;
      RECT 4.240000 1.755000 4.530000 1.800000 ;
      RECT 4.240000 1.940000 4.530000 1.985000 ;
      RECT 4.675000 1.415000 4.965000 1.460000 ;
      RECT 4.675000 1.600000 4.965000 1.645000 ;
  END
END sky130_fd_sc_hd__dfxbp_2
MACRO sky130_fd_sc_hd__dfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.370000 0.715000 1.650000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.890000 1.495000 7.300000 1.575000 ;
        RECT 6.890000 1.575000 7.220000 2.420000 ;
        RECT 6.900000 0.305000 7.230000 0.740000 ;
        RECT 6.900000 0.740000 7.300000 0.825000 ;
        RECT 7.055000 0.825000 7.300000 0.865000 ;
        RECT 7.065000 1.445000 7.300000 1.495000 ;
        RECT 7.110000 0.865000 7.300000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.315000 1.480000 8.650000 2.465000 ;
        RECT 8.395000 0.255000 8.650000 0.910000 ;
        RECT 8.415000 0.910000 8.650000 1.480000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.840000 0.805000 ;
      RECT 0.175000  1.795000 0.840000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.840000 1.795000 ;
      RECT 1.015000  0.345000 1.200000 2.465000 ;
      RECT 1.440000  2.175000 1.705000 2.635000 ;
      RECT 1.455000  0.085000 1.705000 0.545000 ;
      RECT 1.820000  0.675000 2.045000 0.805000 ;
      RECT 1.820000  0.805000 1.990000 1.910000 ;
      RECT 1.820000  1.910000 2.125000 2.040000 ;
      RECT 1.875000  0.365000 2.210000 0.535000 ;
      RECT 1.875000  0.535000 2.045000 0.675000 ;
      RECT 1.875000  2.040000 2.125000 2.465000 ;
      RECT 2.160000  1.125000 2.400000 1.720000 ;
      RECT 2.215000  0.735000 2.740000 0.955000 ;
      RECT 2.335000  2.190000 3.440000 2.360000 ;
      RECT 2.405000  0.365000 3.080000 0.535000 ;
      RECT 2.570000  0.955000 2.740000 1.655000 ;
      RECT 2.570000  1.655000 3.100000 2.020000 ;
      RECT 2.910000  0.535000 3.080000 1.315000 ;
      RECT 2.910000  1.315000 3.780000 1.485000 ;
      RECT 3.270000  1.485000 3.780000 1.575000 ;
      RECT 3.270000  1.575000 3.440000 2.190000 ;
      RECT 3.290000  0.765000 4.120000 1.065000 ;
      RECT 3.290000  1.065000 3.490000 1.095000 ;
      RECT 3.400000  0.085000 3.770000 0.585000 ;
      RECT 3.610000  1.245000 3.780000 1.315000 ;
      RECT 3.610000  1.835000 3.780000 2.635000 ;
      RECT 3.950000  0.365000 4.355000 0.535000 ;
      RECT 3.950000  0.535000 4.120000 0.765000 ;
      RECT 3.950000  1.065000 4.120000 2.135000 ;
      RECT 3.950000  2.135000 4.200000 2.465000 ;
      RECT 4.290000  1.245000 4.480000 1.965000 ;
      RECT 4.425000  2.165000 5.310000 2.335000 ;
      RECT 4.505000  0.705000 4.970000 1.035000 ;
      RECT 4.525000  0.365000 5.310000 0.535000 ;
      RECT 4.650000  1.035000 4.970000 1.995000 ;
      RECT 5.140000  0.535000 5.310000 0.995000 ;
      RECT 5.140000  0.995000 6.020000 1.325000 ;
      RECT 5.140000  1.325000 5.310000 2.165000 ;
      RECT 5.480000  1.530000 6.380000 1.905000 ;
      RECT 5.490000  2.135000 5.805000 2.635000 ;
      RECT 5.585000  0.085000 5.795000 0.615000 ;
      RECT 6.040000  1.905000 6.380000 2.465000 ;
      RECT 6.060000  0.300000 6.390000 0.825000 ;
      RECT 6.190000  0.825000 6.390000 0.995000 ;
      RECT 6.190000  0.995000 6.940000 1.325000 ;
      RECT 6.190000  1.325000 6.380000 1.530000 ;
      RECT 6.550000  1.625000 6.720000 2.635000 ;
      RECT 6.560000  0.085000 6.730000 0.695000 ;
      RECT 7.410000  1.715000 7.740000 2.445000 ;
      RECT 7.420000  0.345000 7.670000 0.615000 ;
      RECT 7.470000  0.615000 7.670000 0.995000 ;
      RECT 7.470000  0.995000 8.245000 1.325000 ;
      RECT 7.470000  1.325000 7.740000 1.715000 ;
      RECT 7.905000  0.085000 8.225000 0.545000 ;
      RECT 7.930000  1.495000 8.145000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.630000  1.785000 0.800000 1.955000 ;
      RECT 1.025000  1.445000 1.195000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.215000  1.445000 2.385000 1.615000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.730000  1.785000 2.900000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.300000  1.785000 4.470000 1.955000 ;
      RECT 4.735000  1.445000 4.905000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
    LAYER met1 ;
      RECT 0.570000 1.755000 0.860000 1.800000 ;
      RECT 0.570000 1.800000 4.530000 1.940000 ;
      RECT 0.570000 1.940000 0.860000 1.985000 ;
      RECT 0.965000 1.415000 1.255000 1.460000 ;
      RECT 0.965000 1.460000 4.965000 1.600000 ;
      RECT 0.965000 1.600000 1.255000 1.645000 ;
      RECT 2.155000 1.415000 2.445000 1.460000 ;
      RECT 2.155000 1.600000 2.445000 1.645000 ;
      RECT 2.670000 1.755000 2.960000 1.800000 ;
      RECT 2.670000 1.940000 2.960000 1.985000 ;
      RECT 4.240000 1.755000 4.530000 1.800000 ;
      RECT 4.240000 1.940000 4.530000 1.985000 ;
      RECT 4.675000 1.415000 4.965000 1.460000 ;
      RECT 4.675000 1.600000 4.965000 1.645000 ;
  END
END sky130_fd_sc_hd__dfxbp_1
MACRO sky130_fd_sc_hd__clkdlybuf4s15_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s15_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.560000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.376300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.210000 0.285000 3.595000 0.545000 ;
        RECT 3.210000 1.760000 3.595000 2.465000 ;
        RECT 3.365000 0.545000 3.595000 1.760000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.255000 0.425000 0.715000 ;
      RECT 0.085000  0.715000 1.215000 0.885000 ;
      RECT 0.085000  1.495000 1.215000 1.665000 ;
      RECT 0.085000  1.665000 0.425000 2.465000 ;
      RECT 0.595000  0.085000 0.910000 0.545000 ;
      RECT 0.595000  1.835000 0.925000 2.635000 ;
      RECT 0.730000  0.885000 1.215000 1.495000 ;
      RECT 1.385000  0.255000 1.760000 0.825000 ;
      RECT 1.385000  1.835000 1.760000 2.465000 ;
      RECT 1.590000  0.825000 1.760000 1.055000 ;
      RECT 1.590000  1.055000 2.685000 1.250000 ;
      RECT 1.590000  1.250000 1.760000 1.835000 ;
      RECT 1.930000  0.255000 2.260000 0.715000 ;
      RECT 1.930000  0.715000 3.195000 0.885000 ;
      RECT 1.930000  1.420000 3.195000 1.590000 ;
      RECT 1.930000  1.590000 2.410000 2.465000 ;
      RECT 2.640000  1.760000 3.040000 2.635000 ;
      RECT 2.710000  0.085000 3.040000 0.545000 ;
      RECT 2.855000  0.885000 3.195000 1.420000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s15_1
MACRO sky130_fd_sc_hd__clkdlybuf4s15_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s15_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.060000 0.555000 1.625000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.397600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.050000 0.255000 3.550000 0.640000 ;
        RECT 3.070000 1.485000 3.550000 2.465000 ;
        RECT 3.355000 0.640000 3.550000 1.485000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.255000 0.415000 0.720000 ;
      RECT 0.085000  0.720000 1.060000 0.890000 ;
      RECT 0.085000  1.795000 1.060000 1.965000 ;
      RECT 0.085000  1.965000 0.430000 2.465000 ;
      RECT 0.585000  0.085000 0.915000 0.550000 ;
      RECT 0.600000  2.135000 0.930000 2.635000 ;
      RECT 0.890000  0.890000 1.060000 1.075000 ;
      RECT 0.890000  1.075000 1.320000 1.245000 ;
      RECT 0.890000  1.245000 1.060000 1.795000 ;
      RECT 1.230000  1.785000 1.660000 2.465000 ;
      RECT 1.280000  0.255000 1.660000 0.905000 ;
      RECT 1.490000  0.905000 1.660000 1.075000 ;
      RECT 1.490000  1.075000 2.415000 1.485000 ;
      RECT 1.490000  1.485000 1.660000 1.785000 ;
      RECT 1.830000  0.255000 2.100000 0.735000 ;
      RECT 1.830000  0.735000 2.900000 0.905000 ;
      RECT 1.830000  1.790000 2.900000 1.965000 ;
      RECT 1.830000  1.965000 2.100000 2.465000 ;
      RECT 2.550000  0.085000 2.880000 0.565000 ;
      RECT 2.550000  2.135000 2.880000 2.635000 ;
      RECT 2.730000  0.905000 2.900000 1.075000 ;
      RECT 2.730000  1.075000 3.185000 1.245000 ;
      RECT 2.730000  1.245000 2.900000 1.790000 ;
      RECT 3.720000  0.085000 4.055000 0.645000 ;
      RECT 3.720000  1.485000 4.055000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s15_2
MACRO sky130_fd_sc_hd__a41o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.785000 0.730000 4.005000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.085000 1.075000 3.550000 1.245000 ;
        RECT 3.335000 0.745000 3.550000 1.075000 ;
        RECT 3.335000 1.245000 3.550000 1.625000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685000 0.995000 2.855000 1.435000 ;
        RECT 2.685000 1.435000 3.090000 1.625000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.000000 0.995000 2.335000 1.625000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.400000 1.075000 1.730000 1.295000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.295000 0.765000 0.755000 ;
        RECT 0.595000 0.755000 0.785000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.805000 ;
      RECT 0.095000  1.495000 0.425000 2.635000 ;
      RECT 0.935000  0.085000 1.265000 0.465000 ;
      RECT 0.980000  0.635000 2.545000 0.805000 ;
      RECT 0.980000  0.805000 1.150000 1.495000 ;
      RECT 0.980000  1.495000 1.785000 1.665000 ;
      RECT 1.015000  1.835000 1.265000 2.635000 ;
      RECT 1.455000  1.665000 1.785000 2.425000 ;
      RECT 1.495000  0.255000 1.705000 0.635000 ;
      RECT 1.875000  0.085000 2.205000 0.465000 ;
      RECT 1.955000  1.795000 3.965000 1.965000 ;
      RECT 1.955000  1.965000 2.125000 2.465000 ;
      RECT 2.335000  2.175000 2.585000 2.635000 ;
      RECT 2.375000  0.295000 4.045000 0.465000 ;
      RECT 2.375000  0.465000 2.545000 0.635000 ;
      RECT 2.795000  1.965000 2.965000 2.465000 ;
      RECT 3.335000  2.175000 3.585000 2.635000 ;
      RECT 3.795000  1.965000 3.965000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a41o_2
MACRO sky130_fd_sc_hd__a41o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 1.075000 4.065000 1.295000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.275000 1.075000 4.975000 1.285000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.155000 1.075000 6.185000 1.295000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.495000 1.075000 7.505000 1.295000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.135000 1.075000 3.145000 1.280000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.635000 1.605000 0.805000 ;
        RECT 0.150000 0.805000 0.320000 1.575000 ;
        RECT 0.150000 1.575000 1.605000 1.745000 ;
        RECT 0.595000 0.255000 0.765000 0.635000 ;
        RECT 0.595000 1.745000 0.765000 2.465000 ;
        RECT 1.435000 0.255000 1.605000 0.635000 ;
        RECT 1.435000 1.745000 1.605000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.095000  1.915000 0.425000 2.635000 ;
      RECT 0.490000  1.075000 1.945000 1.245000 ;
      RECT 0.935000  0.085000 1.265000 0.465000 ;
      RECT 0.935000  1.915000 1.265000 2.635000 ;
      RECT 1.775000  0.085000 2.125000 0.465000 ;
      RECT 1.775000  0.645000 3.905000 0.815000 ;
      RECT 1.775000  0.815000 1.945000 1.075000 ;
      RECT 1.775000  1.245000 1.945000 1.455000 ;
      RECT 1.775000  1.455000 2.965000 1.625000 ;
      RECT 1.775000  1.915000 2.125000 2.635000 ;
      RECT 2.295000  0.255000 2.465000 0.645000 ;
      RECT 2.375000  1.795000 2.545000 2.295000 ;
      RECT 2.375000  2.295000 3.405000 2.465000 ;
      RECT 2.635000  0.085000 2.965000 0.465000 ;
      RECT 2.715000  1.955000 3.045000 2.125000 ;
      RECT 2.795000  1.625000 2.965000 1.955000 ;
      RECT 3.155000  0.295000 4.245000 0.465000 ;
      RECT 3.235000  1.535000 7.370000 1.705000 ;
      RECT 3.235000  1.705000 3.405000 2.295000 ;
      RECT 3.575000  1.915000 3.905000 2.635000 ;
      RECT 4.075000  0.465000 4.245000 0.645000 ;
      RECT 4.075000  0.645000 5.165000 0.815000 ;
      RECT 4.075000  1.705000 4.245000 2.465000 ;
      RECT 4.415000  0.295000 6.105000 0.465000 ;
      RECT 4.415000  1.915000 4.745000 2.635000 ;
      RECT 4.935000  1.705000 5.105000 2.465000 ;
      RECT 5.345000  1.915000 6.035000 2.635000 ;
      RECT 5.355000  0.645000 7.285000 0.815000 ;
      RECT 6.275000  1.705000 6.445000 2.465000 ;
      RECT 6.615000  0.085000 6.945000 0.465000 ;
      RECT 6.615000  1.915000 6.945000 2.635000 ;
      RECT 7.115000  0.255000 7.285000 0.645000 ;
      RECT 7.115000  1.705000 7.285000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__a41o_4
MACRO sky130_fd_sc_hd__a41o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 0.995000 1.915000 1.325000 ;
        RECT 1.535000 1.325000 1.835000 1.620000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.700000 0.415000 2.650000 0.600000 ;
        RECT 2.225000 0.600000 2.445000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705000 0.995000 3.085000 1.625000 ;
        RECT 2.880000 0.395000 3.085000 0.995000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 0.995000 3.570000 1.625000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.075000 1.335000 1.635000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.300000 0.425000 0.560000 ;
        RECT 0.085000 0.560000 0.345000 2.165000 ;
        RECT 0.085000 2.165000 0.425000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.515000  0.735000 1.530000 0.810000 ;
      RECT 0.515000  0.810000 1.335000 0.905000 ;
      RECT 0.515000  0.905000 0.685000 1.825000 ;
      RECT 0.515000  1.825000 1.365000 1.995000 ;
      RECT 0.595000  0.085000 0.925000 0.565000 ;
      RECT 0.595000  2.175000 0.845000 2.635000 ;
      RECT 1.035000  1.995000 1.365000 2.425000 ;
      RECT 1.115000  0.300000 1.530000 0.735000 ;
      RECT 1.535000  1.795000 3.505000 1.965000 ;
      RECT 1.535000  1.965000 1.705000 2.465000 ;
      RECT 1.915000  2.175000 2.165000 2.635000 ;
      RECT 2.375000  1.965000 2.545000 2.465000 ;
      RECT 2.845000  2.175000 3.095000 2.635000 ;
      RECT 3.255000  0.085000 3.595000 0.810000 ;
      RECT 3.335000  1.965000 3.505000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a41o_1
MACRO sky130_fd_sc_hd__o2111ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.820000 1.075000 9.575000 1.340000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.110000 1.075000 7.325000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 1.075000 5.455000 1.345000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 1.075000 3.550000 1.345000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.075000 1.755000 1.345000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  2.984350 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.645000 1.685000 0.815000 ;
        RECT 0.085000 0.815000 0.375000 1.515000 ;
        RECT 0.085000 1.515000 7.390000 1.685000 ;
        RECT 0.085000 1.685000 0.360000 2.465000 ;
        RECT 1.015000 1.685000 1.195000 2.465000 ;
        RECT 1.845000 1.685000 2.035000 2.465000 ;
        RECT 2.685000 1.685000 2.875000 2.465000 ;
        RECT 3.525000 1.685000 3.715000 2.465000 ;
        RECT 4.570000 1.685000 4.760000 2.465000 ;
        RECT 5.410000 1.685000 5.600000 2.465000 ;
        RECT 6.285000 1.685000 6.480000 2.100000 ;
        RECT 7.045000 1.685000 7.390000 1.720000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.095000  0.285000 2.025000 0.475000 ;
      RECT 0.530000  1.855000 0.845000 2.635000 ;
      RECT 1.390000  1.855000 1.675000 2.635000 ;
      RECT 1.855000  0.475000 2.025000 0.615000 ;
      RECT 1.855000  0.615000 3.785000 0.825000 ;
      RECT 2.195000  0.255000 5.565000 0.445000 ;
      RECT 2.205000  1.855000 2.515000 2.635000 ;
      RECT 3.045000  1.855000 3.355000 2.635000 ;
      RECT 3.975000  0.655000 9.440000 0.905000 ;
      RECT 4.075000  1.855000 4.400000 2.635000 ;
      RECT 4.930000  1.855000 5.220000 2.635000 ;
      RECT 5.785000  1.855000 6.115000 2.270000 ;
      RECT 5.785000  2.270000 7.005000 2.465000 ;
      RECT 6.100000  0.085000 6.430000 0.485000 ;
      RECT 6.705000  1.890000 8.235000 2.060000 ;
      RECT 6.705000  2.060000 7.005000 2.270000 ;
      RECT 6.960000  0.085000 7.290000 0.485000 ;
      RECT 7.555000  2.230000 7.885000 2.635000 ;
      RECT 7.825000  0.085000 8.155000 0.485000 ;
      RECT 8.045000  1.515000 9.080000 1.685000 ;
      RECT 8.045000  1.685000 8.235000 1.890000 ;
      RECT 8.055000  2.060000 8.235000 2.465000 ;
      RECT 8.410000  1.855000 8.720000 2.635000 ;
      RECT 8.665000  0.085000 8.995000 0.485000 ;
      RECT 8.890000  1.685000 9.080000 2.465000 ;
      RECT 9.265000  1.535000 9.575000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__o2111ai_4
MACRO sky130_fd_sc_hd__o2111ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 1.005000 3.115000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.995000 2.615000 1.615000 ;
        RECT 2.270000 1.615000 2.615000 2.370000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 1.815000 1.615000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 0.255000 1.355000 1.615000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485000 1.075000 0.815000 1.615000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  0.857250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.690000 0.885000 ;
        RECT 0.085000 0.885000 0.315000 1.785000 ;
        RECT 0.085000 1.785000 2.095000 2.025000 ;
        RECT 0.790000 2.025000 1.025000 2.465000 ;
        RECT 1.750000 2.025000 2.095000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.290000  2.195000 0.620000 2.635000 ;
      RECT 1.210000  2.255000 1.540000 2.635000 ;
      RECT 1.750000  0.255000 2.095000 0.625000 ;
      RECT 1.750000  0.625000 3.115000 0.825000 ;
      RECT 2.285000  0.085000 2.615000 0.455000 ;
      RECT 2.785000  0.255000 3.115000 0.625000 ;
      RECT 2.785000  1.795000 3.115000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o2111ai_1
MACRO sky130_fd_sc_hd__o2111ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635000 1.075000 5.435000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.075000 4.455000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.200000 1.075000 3.185000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.075000 1.790000 1.325000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.355000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.302000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.615000 0.935000 0.905000 ;
        RECT 0.605000 0.905000 0.865000 1.495000 ;
        RECT 0.605000 1.495000 4.005000 1.665000 ;
        RECT 0.605000 1.665000 0.865000 2.465000 ;
        RECT 1.535000 1.665000 1.725000 2.465000 ;
        RECT 2.395000 1.665000 2.575000 2.465000 ;
        RECT 3.815000 1.665000 4.005000 2.105000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.175000  0.260000 1.300000 0.445000 ;
      RECT 0.175000  0.445000 0.435000 0.865000 ;
      RECT 0.175000  1.525000 0.425000 2.635000 ;
      RECT 1.035000  1.835000 1.365000 2.635000 ;
      RECT 1.115000  0.445000 1.300000 0.735000 ;
      RECT 1.115000  0.735000 2.275000 0.905000 ;
      RECT 1.470000  0.255000 3.210000 0.445000 ;
      RECT 1.470000  0.445000 1.775000 0.530000 ;
      RECT 1.470000  0.530000 1.760000 0.565000 ;
      RECT 1.895000  1.840000 2.225000 2.635000 ;
      RECT 1.925000  0.620000 2.275000 0.735000 ;
      RECT 2.450000  0.655000 5.435000 0.840000 ;
      RECT 2.755000  1.835000 3.085000 2.635000 ;
      RECT 2.880000  0.445000 3.210000 0.485000 ;
      RECT 3.310000  1.835000 3.570000 2.275000 ;
      RECT 3.310000  2.275000 4.500000 2.465000 ;
      RECT 3.380000  0.365000 3.570000 0.655000 ;
      RECT 3.740000  0.085000 4.070000 0.485000 ;
      RECT 4.240000  0.365000 4.430000 0.650000 ;
      RECT 4.240000  0.650000 5.435000 0.655000 ;
      RECT 4.240000  1.515000 5.360000 1.685000 ;
      RECT 4.240000  1.685000 4.500000 2.275000 ;
      RECT 4.600000  0.085000 4.930000 0.480000 ;
      RECT 4.670000  1.855000 4.930000 2.635000 ;
      RECT 5.100000  0.365000 5.435000 0.650000 ;
      RECT 5.100000  1.685000 5.360000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__o2111ai_2
MACRO sky130_fd_sc_hd__dlymetal6s4s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s4s_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.570000 1.700000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.660000 0.255000 3.105000 0.825000 ;
        RECT 2.660000 1.495000 3.565000 1.675000 ;
        RECT 2.660000 1.675000 3.105000 2.465000 ;
        RECT 2.735000 0.825000 3.105000 0.995000 ;
        RECT 2.735000 0.995000 3.565000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120000 -0.085000 0.290000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.255000 0.520000 0.655000 ;
      RECT 0.085000  0.655000 1.075000 0.825000 ;
      RECT 0.085000  1.870000 1.075000 2.040000 ;
      RECT 0.085000  2.040000 0.520000 2.465000 ;
      RECT 0.690000  0.085000 1.075000 0.485000 ;
      RECT 0.690000  2.210000 1.075000 2.635000 ;
      RECT 0.740000  0.825000 1.075000 0.995000 ;
      RECT 0.740000  0.995000 1.150000 1.325000 ;
      RECT 0.740000  1.325000 1.075000 1.870000 ;
      RECT 1.245000  0.255000 1.515000 0.825000 ;
      RECT 1.245000  1.495000 1.970000 1.675000 ;
      RECT 1.245000  1.675000 1.515000 2.465000 ;
      RECT 1.320000  0.825000 1.515000 0.995000 ;
      RECT 1.320000  0.995000 1.970000 1.495000 ;
      RECT 1.685000  0.255000 1.935000 0.655000 ;
      RECT 1.685000  0.655000 2.490000 0.825000 ;
      RECT 1.685000  1.845000 2.490000 2.040000 ;
      RECT 1.685000  2.040000 1.935000 2.465000 ;
      RECT 2.105000  0.085000 2.490000 0.485000 ;
      RECT 2.105000  2.210000 2.490000 2.635000 ;
      RECT 2.140000  0.825000 2.490000 0.995000 ;
      RECT 2.140000  0.995000 2.565000 1.325000 ;
      RECT 2.140000  1.325000 2.490000 1.845000 ;
      RECT 3.275000  0.255000 3.530000 0.655000 ;
      RECT 3.275000  0.655000 4.085000 0.825000 ;
      RECT 3.275000  1.845000 4.085000 2.040000 ;
      RECT 3.275000  2.040000 3.530000 2.465000 ;
      RECT 3.700000  0.085000 4.085000 0.485000 ;
      RECT 3.700000  2.210000 4.085000 2.635000 ;
      RECT 3.735000  0.825000 4.085000 0.995000 ;
      RECT 3.735000  0.995000 4.160000 1.325000 ;
      RECT 3.735000  1.325000 4.085000 1.845000 ;
      RECT 4.255000  0.255000 4.515000 0.825000 ;
      RECT 4.255000  1.495000 4.515000 2.465000 ;
      RECT 4.330000  0.825000 4.515000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__dlymetal6s4s_1
MACRO sky130_fd_sc_hd__clkbuf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.745000 0.785000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.383400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 0.255000 1.245000 0.655000 ;
        RECT 1.040000 0.655000 1.725000 0.825000 ;
        RECT 1.060000 1.855000 1.725000 2.030000 ;
        RECT 1.060000 2.030000 1.245000 2.435000 ;
        RECT 1.385000 0.825000 1.725000 1.855000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 1.215000 1.665000 ;
      RECT 0.085000  1.665000 0.355000 2.435000 ;
      RECT 0.525000  1.855000 0.855000 2.635000 ;
      RECT 0.555000  0.085000 0.830000 0.565000 ;
      RECT 0.965000  0.995000 1.215000 1.495000 ;
      RECT 1.415000  0.085000 1.750000 0.485000 ;
      RECT 1.415000  2.210000 1.750000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__clkbuf_2
MACRO sky130_fd_sc_hd__clkbuf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.196500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.985000 1.275000 1.355000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.345000 0.760000 ;
        RECT 0.085000 0.760000 0.255000 1.560000 ;
        RECT 0.085000 1.560000 0.355000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.425000  1.060000 0.710000 1.390000 ;
      RECT 0.525000  0.085000 0.855000 0.465000 ;
      RECT 0.525000  1.875000 0.855000 2.635000 ;
      RECT 0.540000  0.635000 1.205000 0.805000 ;
      RECT 0.540000  0.805000 0.710000 1.060000 ;
      RECT 0.540000  1.390000 0.710000 1.535000 ;
      RECT 0.540000  1.535000 1.205000 1.705000 ;
      RECT 1.035000  0.255000 1.205000 0.635000 ;
      RECT 1.035000  1.705000 1.205000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__clkbuf_1
MACRO sky130_fd_sc_hd__clkbuf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.755000 0.775000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.795200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.345000 1.305000 0.735000 ;
        RECT 1.010000 0.735000 2.660000 0.905000 ;
        RECT 1.045000 1.835000 2.165000 2.005000 ;
        RECT 1.045000 2.005000 1.305000 2.465000 ;
        RECT 1.905000 0.345000 2.165000 0.735000 ;
        RECT 1.905000 1.415000 2.660000 1.585000 ;
        RECT 1.905000 1.585000 2.165000 1.835000 ;
        RECT 1.905000 2.005000 2.165000 2.465000 ;
        RECT 2.255000 0.905000 2.660000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.255000 0.385000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 1.115000 1.665000 ;
      RECT 0.085000  1.665000 0.395000 2.465000 ;
      RECT 0.555000  0.085000 0.830000 0.565000 ;
      RECT 0.565000  1.835000 0.875000 2.635000 ;
      RECT 0.945000  1.075000 2.085000 1.245000 ;
      RECT 0.945000  1.245000 1.115000 1.495000 ;
      RECT 1.475000  0.085000 1.730000 0.565000 ;
      RECT 1.475000  2.175000 1.730000 2.635000 ;
      RECT 2.335000  0.085000 2.615000 0.565000 ;
      RECT 2.335000  1.765000 2.620000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__clkbuf_4
MACRO sky130_fd_sc_hd__clkbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.852000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.400000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.280000 0.280000 2.540000 0.735000 ;
        RECT 2.280000 0.735000 9.025000 0.905000 ;
        RECT 2.280000 1.495000 9.025000 1.720000 ;
        RECT 2.280000 1.720000 7.685000 1.735000 ;
        RECT 2.280000 1.735000 2.540000 2.460000 ;
        RECT 3.140000 0.280000 3.400000 0.735000 ;
        RECT 3.140000 1.735000 3.400000 2.460000 ;
        RECT 4.000000 0.280000 4.260000 0.735000 ;
        RECT 4.000000 1.735000 4.260000 2.460000 ;
        RECT 4.845000 0.280000 5.120000 0.735000 ;
        RECT 4.860000 1.735000 5.120000 2.460000 ;
        RECT 5.705000 0.280000 5.965000 0.735000 ;
        RECT 5.705000 1.735000 5.965000 2.460000 ;
        RECT 6.565000 0.280000 6.825000 0.735000 ;
        RECT 6.565000 1.735000 6.825000 2.460000 ;
        RECT 7.425000 0.280000 7.685000 0.735000 ;
        RECT 7.425000 1.735000 7.685000 2.460000 ;
        RECT 7.860000 0.905000 9.025000 1.495000 ;
        RECT 8.295000 0.280000 8.555000 0.735000 ;
        RECT 8.295000 1.720000 8.585000 2.460000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.085000  0.085000 0.390000 0.595000 ;
      RECT 0.095000  1.825000 0.390000 2.635000 ;
      RECT 0.570000  0.265000 0.820000 1.075000 ;
      RECT 0.570000  1.075000 7.690000 1.325000 ;
      RECT 0.570000  1.325000 0.815000 2.465000 ;
      RECT 0.990000  0.085000 1.250000 0.610000 ;
      RECT 0.990000  1.825000 1.250000 2.635000 ;
      RECT 1.430000  0.265000 1.680000 1.075000 ;
      RECT 1.430000  1.325000 1.680000 2.460000 ;
      RECT 1.850000  0.085000 2.110000 0.645000 ;
      RECT 1.850000  1.835000 2.110000 2.630000 ;
      RECT 1.850000  2.630000 8.125000 2.635000 ;
      RECT 2.710000  0.085000 2.970000 0.565000 ;
      RECT 2.710000  1.905000 2.970000 2.630000 ;
      RECT 3.570000  0.085000 3.830000 0.565000 ;
      RECT 3.570000  1.905000 3.830000 2.630000 ;
      RECT 4.430000  0.085000 4.675000 0.565000 ;
      RECT 4.430000  1.905000 4.690000 2.630000 ;
      RECT 5.290000  0.085000 5.535000 0.565000 ;
      RECT 5.290000  1.905000 5.535000 2.630000 ;
      RECT 6.145000  0.085000 6.395000 0.565000 ;
      RECT 6.150000  1.905000 6.395000 2.630000 ;
      RECT 7.005000  0.085000 7.255000 0.565000 ;
      RECT 7.010000  1.905000 7.255000 2.630000 ;
      RECT 7.865000  0.085000 8.125000 0.565000 ;
      RECT 7.870000  1.905000 8.125000 2.630000 ;
      RECT 8.725000  0.085000 9.025000 0.565000 ;
      RECT 8.755000  1.890000 9.025000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
END sky130_fd_sc_hd__clkbuf_16
MACRO sky130_fd_sc_hd__clkbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.426000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 0.400000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.590400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 0.280000 1.680000 0.735000 ;
        RECT 1.420000 0.735000 4.730000 0.905000 ;
        RECT 1.420000 1.495000 4.730000 1.735000 ;
        RECT 1.420000 1.735000 1.680000 2.460000 ;
        RECT 2.280000 0.280000 2.540000 0.735000 ;
        RECT 2.280000 1.735000 2.540000 2.460000 ;
        RECT 3.140000 0.280000 3.400000 0.735000 ;
        RECT 3.140000 1.735000 3.400000 2.460000 ;
        RECT 3.760000 0.905000 4.730000 1.495000 ;
        RECT 4.000000 0.280000 4.260000 0.735000 ;
        RECT 4.000000 1.735000 4.260000 2.460000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.095000  1.525000 0.390000 2.635000 ;
      RECT 0.145000  0.085000 0.390000 0.545000 ;
      RECT 0.570000  0.265000 0.820000 1.075000 ;
      RECT 0.570000  1.075000 3.590000 1.325000 ;
      RECT 0.570000  1.325000 0.820000 2.460000 ;
      RECT 0.990000  0.085000 1.250000 0.610000 ;
      RECT 0.990000  1.525000 1.250000 2.635000 ;
      RECT 1.850000  0.085000 2.110000 0.565000 ;
      RECT 1.850000  1.905000 2.110000 2.635000 ;
      RECT 2.710000  0.085000 2.970000 0.565000 ;
      RECT 2.710000  1.905000 2.970000 2.635000 ;
      RECT 3.570000  0.085000 3.830000 0.565000 ;
      RECT 3.570000  1.905000 3.830000 2.635000 ;
      RECT 4.430000  0.085000 4.730000 0.565000 ;
      RECT 4.430000  1.905000 4.725000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__clkbuf_8
MACRO sky130_fd_sc_hd__and3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.635000 0.635000 1.020000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 2.125000 1.345000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.145000 0.305000 1.365000 0.790000 ;
        RECT 1.145000 0.790000 1.475000 1.215000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 1.765000 2.215000 2.465000 ;
        RECT 1.955000 0.255000 2.215000 0.735000 ;
        RECT 2.045000 0.735000 2.215000 1.765000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.295000 0.975000 0.465000 ;
      RECT 0.085000  1.190000 0.975000 1.260000 ;
      RECT 0.085000  1.260000 0.980000 1.285000 ;
      RECT 0.085000  1.285000 0.990000 1.300000 ;
      RECT 0.085000  1.300000 0.995000 1.315000 ;
      RECT 0.085000  1.315000 1.005000 1.320000 ;
      RECT 0.085000  1.320000 1.010000 1.330000 ;
      RECT 0.085000  1.330000 1.015000 1.340000 ;
      RECT 0.085000  1.340000 1.025000 1.345000 ;
      RECT 0.085000  1.345000 1.035000 1.355000 ;
      RECT 0.085000  1.355000 1.045000 1.360000 ;
      RECT 0.085000  1.360000 0.345000 1.810000 ;
      RECT 0.085000  1.980000 0.700000 2.080000 ;
      RECT 0.085000  2.080000 0.690000 2.635000 ;
      RECT 0.515000  1.710000 0.845000 1.955000 ;
      RECT 0.515000  1.955000 0.700000 1.980000 ;
      RECT 0.710000  1.360000 1.045000 1.365000 ;
      RECT 0.710000  1.365000 1.060000 1.370000 ;
      RECT 0.710000  1.370000 1.075000 1.380000 ;
      RECT 0.710000  1.380000 1.100000 1.385000 ;
      RECT 0.710000  1.385000 1.875000 1.390000 ;
      RECT 0.740000  1.390000 1.875000 1.425000 ;
      RECT 0.775000  1.425000 1.875000 1.450000 ;
      RECT 0.805000  0.465000 0.975000 1.190000 ;
      RECT 0.805000  1.450000 1.875000 1.480000 ;
      RECT 0.825000  1.480000 1.875000 1.510000 ;
      RECT 0.845000  1.510000 1.875000 1.540000 ;
      RECT 0.915000  1.540000 1.875000 1.550000 ;
      RECT 0.940000  1.550000 1.875000 1.560000 ;
      RECT 0.960000  1.560000 1.875000 1.575000 ;
      RECT 0.980000  1.575000 1.875000 1.590000 ;
      RECT 0.985000  1.590000 1.770000 1.600000 ;
      RECT 1.000000  1.600000 1.770000 1.635000 ;
      RECT 1.015000  1.635000 1.770000 1.885000 ;
      RECT 1.515000  2.090000 1.770000 2.635000 ;
      RECT 1.535000  0.085000 1.785000 0.625000 ;
      RECT 1.645000  0.990000 1.875000 1.385000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__and3_1
MACRO sky130_fd_sc_hd__and3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.470000 1.245000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.895000 2.125000 1.370000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.305000 1.295000 0.750000 ;
        RECT 1.065000 0.750000 1.475000 1.245000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 1.795000 2.245000 2.465000 ;
        RECT 1.980000 0.255000 2.230000 0.715000 ;
        RECT 2.060000 0.715000 2.230000 0.925000 ;
        RECT 2.060000 0.925000 2.675000 1.445000 ;
        RECT 2.075000 1.445000 2.245000 1.795000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  2.130000 0.715000 2.635000 ;
      RECT 0.100000  1.425000 1.890000 1.595000 ;
      RECT 0.100000  1.595000 0.355000 1.960000 ;
      RECT 0.105000  0.305000 0.895000 0.570000 ;
      RECT 0.525000  1.765000 0.855000 1.955000 ;
      RECT 0.525000  1.955000 0.715000 2.130000 ;
      RECT 0.640000  0.570000 0.895000 1.425000 ;
      RECT 1.080000  1.595000 1.330000 1.890000 ;
      RECT 1.475000  0.085000 1.805000 0.580000 ;
      RECT 1.555000  1.790000 1.770000 2.635000 ;
      RECT 1.660000  0.995000 1.890000 1.425000 ;
      RECT 2.400000  0.085000 2.675000 0.745000 ;
      RECT 2.415000  1.625000 2.675000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__and3_2
MACRO sky130_fd_sc_hd__and3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.995000 0.875000 1.340000 ;
        RECT 0.115000 1.340000 0.365000 2.335000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.745000 1.355000 1.340000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 1.900000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.450000 0.515000 2.640000 0.615000 ;
        RECT 2.450000 0.615000 4.055000 0.845000 ;
        RECT 2.450000 1.535000 4.055000 1.760000 ;
        RECT 2.450000 1.760000 2.640000 2.465000 ;
        RECT 3.310000 0.255000 3.500000 0.615000 ;
        RECT 3.310000 1.760000 4.055000 1.765000 ;
        RECT 3.310000 1.765000 3.500000 2.465000 ;
        RECT 3.775000 0.845000 4.055000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.465000  0.255000 0.800000 0.375000 ;
      RECT 0.465000  0.375000 1.725000 0.565000 ;
      RECT 0.465000  0.565000 0.800000 0.805000 ;
      RECT 0.545000  1.580000 2.280000 1.750000 ;
      RECT 0.545000  1.750000 0.725000 2.465000 ;
      RECT 0.895000  1.935000 1.345000 2.635000 ;
      RECT 1.520000  1.750000 1.700000 2.465000 ;
      RECT 1.535000  0.565000 1.725000 0.615000 ;
      RECT 1.535000  0.615000 2.280000 0.805000 ;
      RECT 1.905000  0.085000 2.235000 0.445000 ;
      RECT 1.910000  1.935000 2.240000 2.635000 ;
      RECT 2.070000  0.805000 2.280000 1.020000 ;
      RECT 2.070000  1.020000 3.605000 1.355000 ;
      RECT 2.070000  1.355000 2.280000 1.580000 ;
      RECT 2.810000  0.085000 3.140000 0.445000 ;
      RECT 2.810000  1.935000 3.140000 2.635000 ;
      RECT 3.670000  0.085000 4.000000 0.445000 ;
      RECT 3.670000  1.935000 4.000000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__and3_4
MACRO sky130_fd_sc_hd__diode_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__diode_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.920000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIODE
    ANTENNADIFFAREA  0.434700 ;
    ANTENNAGATEAREA  0.434700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.835000 2.465000 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.920000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.110000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.920000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.920000 0.085000 ;
      RECT 0.000000  2.635000 0.920000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
  END
END sky130_fd_sc_hd__diode_2
MACRO sky130_fd_sc_hd__a31o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 0.995000 2.160000 1.655000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 0.995000 1.700000 1.655000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 0.995000 1.240000 1.325000 ;
        RECT 1.025000 1.325000 1.240000 1.655000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 0.995000 2.620000 1.655000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.437250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.300000 0.425000 0.810000 ;
        RECT 0.095000 0.810000 0.285000 1.575000 ;
        RECT 0.095000 1.575000 0.425000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.455000  0.995000 0.765000 1.325000 ;
      RECT 0.595000  0.085000 0.925000 0.485000 ;
      RECT 0.595000  0.655000 2.960000 0.825000 ;
      RECT 0.595000  0.825000 0.765000 0.995000 ;
      RECT 0.595000  1.495000 0.845000 2.635000 ;
      RECT 1.035000  1.825000 2.325000 1.995000 ;
      RECT 1.035000  1.995000 1.285000 2.415000 ;
      RECT 1.515000  2.165000 1.845000 2.635000 ;
      RECT 1.975000  0.315000 2.305000 0.655000 ;
      RECT 2.075000  1.995000 2.325000 2.415000 ;
      RECT 2.475000  0.085000 2.805000 0.485000 ;
      RECT 2.505000  1.825000 2.960000 1.995000 ;
      RECT 2.505000  1.995000 2.835000 2.425000 ;
      RECT 2.790000  0.825000 2.960000 1.825000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a31o_1
MACRO sky130_fd_sc_hd__a31o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 0.415000 2.175000 0.700000 ;
        RECT 1.965000 0.700000 2.355000 0.870000 ;
        RECT 2.185000 0.870000 2.355000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.400000 1.700000 0.695000 ;
        RECT 1.530000 0.695000 1.795000 0.865000 ;
        RECT 1.625000 0.865000 1.795000 1.075000 ;
        RECT 1.625000 1.075000 1.955000 1.245000 ;
        RECT 1.625000 1.245000 1.795000 1.260000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.760000 1.270000 0.995000 ;
        RECT 1.065000 0.995000 1.395000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895000 0.755000 3.090000 1.325000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.715000 0.765000 0.885000 ;
        RECT 0.090000 0.885000 0.345000 1.835000 ;
        RECT 0.090000 1.835000 0.765000 2.005000 ;
        RECT 0.595000 0.255000 0.765000 0.715000 ;
        RECT 0.595000 2.005000 0.765000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.545000 ;
      RECT 0.135000  2.175000 0.385000 2.635000 ;
      RECT 0.555000  1.075000 0.885000 1.245000 ;
      RECT 0.555000  1.245000 0.725000 1.495000 ;
      RECT 0.555000  1.495000 3.045000 1.665000 ;
      RECT 0.935000  1.835000 1.185000 2.635000 ;
      RECT 0.955000  0.085000 1.285000 0.465000 ;
      RECT 1.015000  0.465000 1.185000 0.545000 ;
      RECT 1.355000  1.835000 2.645000 2.005000 ;
      RECT 1.355000  2.005000 1.605000 2.425000 ;
      RECT 1.815000  2.175000 2.145000 2.635000 ;
      RECT 2.335000  2.005000 2.585000 2.425000 ;
      RECT 2.375000  0.335000 2.705000 0.505000 ;
      RECT 2.460000  0.255000 2.705000 0.335000 ;
      RECT 2.535000  0.505000 2.705000 1.495000 ;
      RECT 2.875000  0.085000 3.135000 0.565000 ;
      RECT 2.875000  1.665000 3.045000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a31o_2
MACRO sky130_fd_sc_hd__a31o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.075000 1.705000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.725000 1.075000 1.055000 1.245000 ;
        RECT 0.805000 0.735000 2.170000 0.905000 ;
        RECT 0.805000 0.905000 0.975000 1.075000 ;
        RECT 1.985000 0.905000 2.170000 1.075000 ;
        RECT 1.985000 1.075000 2.315000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 1.075000 0.525000 1.445000 ;
        RECT 0.150000 1.445000 2.855000 1.615000 ;
        RECT 2.525000 1.075000 2.855000 1.445000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.575000 1.075000 4.030000 1.285000 ;
        RECT 3.815000 0.745000 4.030000 1.075000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505000 0.655000 6.295000 0.825000 ;
        RECT 4.535000 1.785000 6.295000 1.955000 ;
        RECT 4.595000 1.955000 4.765000 2.465000 ;
        RECT 5.435000 1.955000 5.605000 2.465000 ;
        RECT 6.125000 0.825000 6.295000 1.785000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.085000 0.345000 0.905000 ;
      RECT 0.175000  1.785000 2.985000 1.955000 ;
      RECT 0.175000  1.955000 0.345000 2.465000 ;
      RECT 0.515000  2.125000 0.845000 2.635000 ;
      RECT 1.015000  1.955000 1.185000 2.465000 ;
      RECT 1.355000  0.395000 2.520000 0.565000 ;
      RECT 1.355000  2.125000 1.685000 2.635000 ;
      RECT 1.855000  1.955000 2.025000 2.465000 ;
      RECT 2.195000  2.125000 2.525000 2.635000 ;
      RECT 2.350000  0.565000 2.520000 0.700000 ;
      RECT 2.350000  0.700000 3.485000 0.805000 ;
      RECT 2.350000  0.805000 3.345000 0.870000 ;
      RECT 2.700000  0.085000 2.985000 0.530000 ;
      RECT 2.815000  1.955000 2.985000 2.295000 ;
      RECT 2.815000  2.295000 3.825000 2.465000 ;
      RECT 3.155000  0.295000 3.485000 0.700000 ;
      RECT 3.155000  0.870000 3.345000 1.455000 ;
      RECT 3.155000  1.455000 4.395000 1.625000 ;
      RECT 3.155000  1.625000 3.485000 2.115000 ;
      RECT 3.655000  1.795000 3.825000 2.295000 ;
      RECT 3.735000  0.085000 4.265000 0.565000 ;
      RECT 4.095000  2.125000 4.425000 2.635000 ;
      RECT 4.225000  0.995000 5.935000 1.325000 ;
      RECT 4.225000  1.325000 4.395000 1.455000 ;
      RECT 4.935000  0.085000 5.265000 0.485000 ;
      RECT 4.935000  2.125000 5.265000 2.635000 ;
      RECT 5.775000  0.085000 6.105000 0.485000 ;
      RECT 5.775000  2.125000 6.105000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__a31o_4
MACRO sky130_fd_sc_hd__sdfbbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfbbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.26000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775000 1.405000 4.105000 1.575000 ;
        RECT 3.775000 1.575000 4.060000 1.675000 ;
        RECT 3.825000 1.675000 4.060000 2.375000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.915000 0.255000 14.175000 0.785000 ;
        RECT 13.915000 1.470000 14.175000 2.465000 ;
        RECT 13.965000 0.785000 14.175000 1.470000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.500000 0.255000 12.785000 0.715000 ;
        RECT 12.500000 1.630000 12.785000 2.465000 ;
        RECT 12.605000 0.715000 12.785000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.535000 1.095000 11.990000 1.325000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 1.025000 1.695000 1.685000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.345000 2.155000 0.815000 ;
        RECT 1.935000 0.815000 2.315000 1.150000 ;
        RECT 1.935000 1.150000 2.155000 1.695000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.870000 0.735000 6.295000 0.965000 ;
        RECT 5.870000 0.965000 6.215000 1.065000 ;
      LAYER mcon ;
        RECT 6.125000 0.765000 6.295000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755000 0.735000 10.130000 1.065000 ;
      LAYER mcon ;
        RECT 9.805000 0.765000 9.975000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065000 0.735000  6.355000 0.780000 ;
        RECT 6.065000 0.780000 10.035000 0.920000 ;
        RECT 6.065000 0.920000  6.355000 0.965000 ;
        RECT 9.745000 0.735000 10.035000 0.780000 ;
        RECT 9.745000 0.920000 10.035000 0.965000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 14.450000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.095000  0.345000  0.345000 0.635000 ;
      RECT  0.095000  0.635000  0.835000 0.805000 ;
      RECT  0.095000  1.795000  0.835000 1.965000 ;
      RECT  0.095000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.605000  0.805000  0.835000 1.795000 ;
      RECT  1.015000  0.345000  1.235000 2.465000 ;
      RECT  1.430000  0.085000  1.705000 0.635000 ;
      RECT  1.430000  1.885000  1.785000 2.635000 ;
      RECT  2.215000  1.875000  2.575000 2.385000 ;
      RECT  2.325000  0.265000  2.655000 0.595000 ;
      RECT  2.405000  1.295000  3.075000 1.405000 ;
      RECT  2.405000  1.405000  2.670000 1.430000 ;
      RECT  2.405000  1.430000  2.630000 1.465000 ;
      RECT  2.405000  1.465000  2.605000 1.505000 ;
      RECT  2.405000  1.505000  2.575000 1.875000 ;
      RECT  2.460000  1.255000  3.075000 1.295000 ;
      RECT  2.485000  0.595000  2.655000 1.075000 ;
      RECT  2.485000  1.075000  3.075000 1.255000 ;
      RECT  2.760000  1.575000  3.605000 1.745000 ;
      RECT  2.760000  1.745000  3.140000 1.905000 ;
      RECT  2.870000  0.305000  3.040000 0.625000 ;
      RECT  2.870000  0.625000  3.645000 0.765000 ;
      RECT  2.870000  0.765000  3.770000 0.795000 ;
      RECT  2.970000  1.905000  3.140000 2.465000 ;
      RECT  3.225000  0.085000  3.555000 0.445000 ;
      RECT  3.310000  2.215000  3.640000 2.635000 ;
      RECT  3.430000  0.795000  3.770000 1.095000 ;
      RECT  3.430000  1.095000  3.605000 1.575000 ;
      RECT  3.950000  0.425000  4.330000 0.595000 ;
      RECT  3.950000  0.595000  4.120000 1.065000 ;
      RECT  3.950000  1.065000  4.400000 1.105000 ;
      RECT  3.950000  1.105000  4.410000 1.175000 ;
      RECT  3.950000  1.175000  4.445000 1.235000 ;
      RECT  4.160000  0.265000  4.330000 0.425000 ;
      RECT  4.225000  1.235000  4.445000 1.275000 ;
      RECT  4.230000  2.135000  4.445000 2.465000 ;
      RECT  4.245000  1.275000  4.445000 1.305000 ;
      RECT  4.275000  1.305000  4.445000 2.135000 ;
      RECT  4.555000  0.265000  5.655000 0.465000 ;
      RECT  4.570000  0.705000  4.790000 1.035000 ;
      RECT  4.615000  1.035000  4.790000 1.575000 ;
      RECT  4.615000  1.575000  5.125000 1.955000 ;
      RECT  4.635000  2.250000  5.465000 2.420000 ;
      RECT  5.000000  0.735000  5.330000 1.015000 ;
      RECT  5.295000  1.195000  5.670000 1.235000 ;
      RECT  5.295000  1.235000  6.645000 1.405000 ;
      RECT  5.295000  1.405000  5.465000 2.250000 ;
      RECT  5.485000  0.465000  5.655000 0.585000 ;
      RECT  5.485000  0.585000  5.670000 0.655000 ;
      RECT  5.500000  0.655000  5.670000 1.195000 ;
      RECT  5.635000  1.575000  5.885000 1.785000 ;
      RECT  5.635000  1.785000  6.985000 2.035000 ;
      RECT  5.705000  2.205000  6.085000 2.635000 ;
      RECT  5.835000  0.085000  6.005000 0.525000 ;
      RECT  6.260000  0.255000  7.350000 0.425000 ;
      RECT  6.260000  0.425000  6.590000 0.465000 ;
      RECT  6.385000  2.035000  6.555000 2.375000 ;
      RECT  6.395000  1.405000  6.645000 1.485000 ;
      RECT  6.425000  1.155000  6.645000 1.235000 ;
      RECT  6.680000  0.610000  7.010000 0.780000 ;
      RECT  6.810000  0.780000  7.010000 0.895000 ;
      RECT  6.810000  0.895000  8.125000 1.060000 ;
      RECT  6.815000  1.060000  8.125000 1.065000 ;
      RECT  6.815000  1.065000  6.985000 1.785000 ;
      RECT  7.155000  1.235000  7.485000 1.415000 ;
      RECT  7.155000  1.415000  8.160000 1.655000 ;
      RECT  7.175000  1.915000  7.505000 2.635000 ;
      RECT  7.180000  0.425000  7.350000 0.715000 ;
      RECT  7.620000  0.085000  7.975000 0.465000 ;
      RECT  7.795000  1.065000  8.125000 1.235000 ;
      RECT  8.360000  1.575000  8.595000 1.985000 ;
      RECT  8.420000  0.705000  8.705000 1.125000 ;
      RECT  8.420000  1.125000  9.040000 1.305000 ;
      RECT  8.550000  2.250000  9.380000 2.420000 ;
      RECT  8.615000  0.265000  9.380000 0.465000 ;
      RECT  8.835000  1.305000  9.040000 1.905000 ;
      RECT  9.210000  0.465000  9.380000 1.235000 ;
      RECT  9.210000  1.235000 10.560000 1.405000 ;
      RECT  9.210000  1.405000  9.380000 2.250000 ;
      RECT  9.550000  1.575000  9.800000 1.915000 ;
      RECT  9.550000  1.915000 12.330000 2.085000 ;
      RECT  9.560000  0.085000  9.820000 0.525000 ;
      RECT  9.620000  2.255000 10.000000 2.635000 ;
      RECT 10.080000  0.255000 11.250000 0.425000 ;
      RECT 10.080000  0.425000 10.410000 0.545000 ;
      RECT 10.240000  2.085000 10.410000 2.375000 ;
      RECT 10.340000  1.075000 10.560000 1.235000 ;
      RECT 10.575000  0.595000 10.905000 0.780000 ;
      RECT 10.730000  0.780000 10.905000 1.915000 ;
      RECT 10.940000  2.255000 12.330000 2.635000 ;
      RECT 11.075000  0.425000 11.250000 0.585000 ;
      RECT 11.080000  0.755000 11.775000 0.925000 ;
      RECT 11.080000  0.925000 11.355000 1.575000 ;
      RECT 11.080000  1.575000 11.855000 1.745000 ;
      RECT 11.565000  0.265000 11.775000 0.755000 ;
      RECT 12.000000  0.085000 12.330000 0.805000 ;
      RECT 12.160000  0.995000 12.425000 1.325000 ;
      RECT 12.160000  1.325000 12.330000 1.915000 ;
      RECT 12.960000  0.255000 13.275000 0.995000 ;
      RECT 12.960000  0.995000 13.795000 1.325000 ;
      RECT 12.960000  1.325000 13.275000 2.415000 ;
      RECT 13.455000  0.085000 13.745000 0.545000 ;
      RECT 13.455000  1.765000 13.740000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  0.765000  0.775000 0.935000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  1.785000  1.235000 1.955000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  1.105000  3.075000 1.275000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.230000  1.105000  4.400000 1.275000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.785000  4.915000 1.955000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.155000  0.765000  5.325000 0.935000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  1.445000  8.135000 1.615000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  1.105000  8.595000 1.275000 ;
      RECT  8.425000  1.785000  8.595000 1.955000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  1.445000 11.355000 1.615000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT  0.545000 0.735000  0.835000 0.780000 ;
      RECT  0.545000 0.780000  5.385000 0.920000 ;
      RECT  0.545000 0.920000  0.835000 0.965000 ;
      RECT  1.005000 1.755000  1.295000 1.800000 ;
      RECT  1.005000 1.800000  8.655000 1.940000 ;
      RECT  1.005000 1.940000  1.295000 1.985000 ;
      RECT  2.845000 1.075000  3.135000 1.120000 ;
      RECT  2.845000 1.120000  4.460000 1.260000 ;
      RECT  2.845000 1.260000  3.135000 1.305000 ;
      RECT  4.170000 1.075000  4.460000 1.120000 ;
      RECT  4.170000 1.260000  4.460000 1.305000 ;
      RECT  4.685000 1.755000  4.975000 1.800000 ;
      RECT  4.685000 1.940000  4.975000 1.985000 ;
      RECT  5.095000 0.735000  5.385000 0.780000 ;
      RECT  5.095000 0.920000  5.385000 0.965000 ;
      RECT  5.170000 0.965000  5.385000 1.120000 ;
      RECT  5.170000 1.120000  8.655000 1.260000 ;
      RECT  7.905000 1.415000  8.195000 1.460000 ;
      RECT  7.905000 1.460000 11.415000 1.600000 ;
      RECT  7.905000 1.600000  8.195000 1.645000 ;
      RECT  8.365000 1.075000  8.655000 1.120000 ;
      RECT  8.365000 1.260000  8.655000 1.305000 ;
      RECT  8.365000 1.755000  8.655000 1.800000 ;
      RECT  8.365000 1.940000  8.655000 1.985000 ;
      RECT 11.125000 1.415000 11.415000 1.460000 ;
      RECT 11.125000 1.600000 11.415000 1.645000 ;
  END
END sky130_fd_sc_hd__sdfbbn_1
MACRO sky130_fd_sc_hd__sdfbbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfbbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.18000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 1.325000 4.025000 2.375000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.415000 0.255000 14.665000 0.825000 ;
        RECT 14.415000 1.445000 14.665000 2.465000 ;
        RECT 14.460000 0.825000 14.665000 1.445000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.580000 0.255000 12.830000 0.715000 ;
        RECT 12.580000 1.630000 12.830000 2.465000 ;
        RECT 12.660000 0.715000 12.830000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.590000 1.095000 12.070000 1.325000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 1.025000 1.695000 1.685000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.345000 2.145000 0.765000 ;
        RECT 1.935000 0.765000 2.335000 1.095000 ;
        RECT 1.935000 1.095000 2.155000 1.695000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 0.735000 6.295000 0.965000 ;
        RECT 5.885000 0.965000 6.215000 1.065000 ;
      LAYER mcon ;
        RECT 6.125000 0.765000 6.295000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755000 0.735000 10.130000 1.065000 ;
      LAYER mcon ;
        RECT 9.805000 0.765000 9.975000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065000 0.735000  6.355000 0.780000 ;
        RECT 6.065000 0.780000 10.035000 0.920000 ;
        RECT 6.065000 0.920000  6.355000 0.965000 ;
        RECT 9.745000 0.735000 10.035000 0.780000 ;
        RECT 9.745000 0.920000 10.035000 0.965000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.180000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 15.370000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 15.180000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.180000 0.085000 ;
      RECT  0.000000  2.635000 15.180000 2.805000 ;
      RECT  0.170000  0.345000  0.345000 0.635000 ;
      RECT  0.170000  0.635000  0.835000 0.805000 ;
      RECT  0.170000  1.795000  0.835000 1.965000 ;
      RECT  0.170000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.605000  0.805000  0.835000 1.795000 ;
      RECT  1.015000  0.345000  1.235000 2.465000 ;
      RECT  1.430000  0.085000  1.705000 0.635000 ;
      RECT  1.430000  1.885000  1.785000 2.635000 ;
      RECT  2.215000  1.875000  2.575000 2.385000 ;
      RECT  2.315000  0.265000  2.730000 0.595000 ;
      RECT  2.405000  1.250000  3.075000 1.405000 ;
      RECT  2.405000  1.405000  2.575000 1.875000 ;
      RECT  2.435000  1.235000  3.075000 1.250000 ;
      RECT  2.560000  0.595000  2.730000 1.075000 ;
      RECT  2.560000  1.075000  3.075000 1.235000 ;
      RECT  2.745000  1.575000  3.645000 1.745000 ;
      RECT  2.745000  1.745000  3.065000 1.905000 ;
      RECT  2.895000  1.905000  3.065000 2.465000 ;
      RECT  2.955000  0.305000  3.125000 0.625000 ;
      RECT  2.955000  0.625000  3.645000 0.765000 ;
      RECT  2.955000  0.765000  3.770000 0.795000 ;
      RECT  3.295000  2.215000  3.640000 2.635000 ;
      RECT  3.370000  0.085000  3.700000 0.445000 ;
      RECT  3.475000  0.795000  3.770000 1.095000 ;
      RECT  3.475000  1.095000  3.645000 1.575000 ;
      RECT  4.230000  0.305000  4.455000 2.465000 ;
      RECT  4.625000  0.705000  4.845000 1.575000 ;
      RECT  4.625000  1.575000  5.125000 1.955000 ;
      RECT  4.635000  2.250000  5.465000 2.420000 ;
      RECT  4.700000  0.265000  5.715000 0.465000 ;
      RECT  5.025000  0.645000  5.375000 1.015000 ;
      RECT  5.295000  1.195000  5.715000 1.235000 ;
      RECT  5.295000  1.235000  6.645000 1.405000 ;
      RECT  5.295000  1.405000  5.465000 2.250000 ;
      RECT  5.545000  0.465000  5.715000 1.195000 ;
      RECT  5.635000  1.575000  5.885000 1.785000 ;
      RECT  5.635000  1.785000  6.985000 2.035000 ;
      RECT  5.705000  2.205000  6.085000 2.635000 ;
      RECT  5.885000  0.085000  6.055000 0.525000 ;
      RECT  6.225000  0.255000  7.375000 0.425000 ;
      RECT  6.225000  0.425000  6.555000 0.505000 ;
      RECT  6.385000  2.035000  6.555000 2.375000 ;
      RECT  6.395000  1.405000  6.645000 1.485000 ;
      RECT  6.425000  1.155000  6.645000 1.235000 ;
      RECT  6.705000  0.595000  7.035000 0.765000 ;
      RECT  6.815000  0.765000  7.035000 0.895000 ;
      RECT  6.815000  0.895000  8.125000 1.065000 ;
      RECT  6.815000  1.065000  6.985000 1.785000 ;
      RECT  7.155000  1.235000  7.485000 1.415000 ;
      RECT  7.155000  1.415000  8.160000 1.655000 ;
      RECT  7.175000  1.915000  7.505000 2.635000 ;
      RECT  7.205000  0.425000  7.375000 0.715000 ;
      RECT  7.645000  0.085000  7.975000 0.465000 ;
      RECT  7.795000  1.065000  8.125000 1.235000 ;
      RECT  8.360000  1.575000  8.595000 1.985000 ;
      RECT  8.420000  0.705000  8.705000 1.125000 ;
      RECT  8.420000  1.125000  9.040000 1.305000 ;
      RECT  8.550000  2.250000  9.380000 2.420000 ;
      RECT  8.615000  0.265000  9.380000 0.465000 ;
      RECT  8.835000  1.305000  9.040000 1.905000 ;
      RECT  9.210000  0.465000  9.380000 1.235000 ;
      RECT  9.210000  1.235000 10.560000 1.405000 ;
      RECT  9.210000  1.405000  9.380000 2.250000 ;
      RECT  9.550000  1.575000  9.800000 1.915000 ;
      RECT  9.550000  1.915000 12.410000 2.085000 ;
      RECT  9.560000  0.085000  9.820000 0.525000 ;
      RECT  9.620000  2.255000 10.000000 2.635000 ;
      RECT 10.080000  0.255000 11.250000 0.425000 ;
      RECT 10.080000  0.425000 10.410000 0.545000 ;
      RECT 10.240000  2.085000 10.410000 2.375000 ;
      RECT 10.340000  1.075000 10.560000 1.235000 ;
      RECT 10.580000  0.595000 10.910000 0.780000 ;
      RECT 10.730000  0.780000 10.910000 1.915000 ;
      RECT 10.940000  2.255000 12.410000 2.635000 ;
      RECT 11.080000  0.425000 11.250000 0.585000 ;
      RECT 11.080000  0.755000 11.845000 0.925000 ;
      RECT 11.080000  0.925000 11.355000 1.575000 ;
      RECT 11.080000  1.575000 11.925000 1.745000 ;
      RECT 11.620000  0.265000 11.845000 0.755000 ;
      RECT 12.080000  0.085000 12.410000 0.805000 ;
      RECT 12.240000  0.995000 12.480000 1.325000 ;
      RECT 12.240000  1.325000 12.410000 1.915000 ;
      RECT 13.000000  0.085000 13.235000 0.885000 ;
      RECT 13.000000  1.495000 13.235000 2.635000 ;
      RECT 13.455000  0.255000 13.770000 0.995000 ;
      RECT 13.455000  0.995000 14.290000 1.325000 ;
      RECT 13.455000  1.325000 13.770000 2.415000 ;
      RECT 13.950000  0.085000 14.245000 0.545000 ;
      RECT 13.950000  1.765000 14.245000 2.635000 ;
      RECT 14.835000  0.085000 15.075000 0.885000 ;
      RECT 14.835000  1.495000 15.075000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  0.765000  0.775000 0.935000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  1.785000  1.235000 1.955000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  1.105000  3.075000 1.275000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.785000  4.915000 1.955000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  0.765000  5.375000 0.935000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  1.445000  8.135000 1.615000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  1.105000  8.595000 1.275000 ;
      RECT  8.425000  1.785000  8.595000 1.955000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  1.445000 11.355000 1.615000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
    LAYER met1 ;
      RECT  0.545000 0.735000  0.835000 0.780000 ;
      RECT  0.545000 0.780000  5.435000 0.920000 ;
      RECT  0.545000 0.920000  0.835000 0.965000 ;
      RECT  1.005000 1.755000  1.295000 1.800000 ;
      RECT  1.005000 1.800000  8.655000 1.940000 ;
      RECT  1.005000 1.940000  1.295000 1.985000 ;
      RECT  2.845000 1.075000  3.135000 1.120000 ;
      RECT  2.845000 1.120000  4.515000 1.260000 ;
      RECT  2.845000 1.260000  3.135000 1.305000 ;
      RECT  4.225000 1.075000  4.515000 1.120000 ;
      RECT  4.225000 1.260000  4.515000 1.305000 ;
      RECT  4.685000 1.755000  4.975000 1.800000 ;
      RECT  4.685000 1.940000  4.975000 1.985000 ;
      RECT  5.145000 0.735000  5.435000 0.780000 ;
      RECT  5.145000 0.920000  5.435000 0.965000 ;
      RECT  5.220000 0.965000  5.435000 1.120000 ;
      RECT  5.220000 1.120000  8.655000 1.260000 ;
      RECT  7.905000 1.415000  8.195000 1.460000 ;
      RECT  7.905000 1.460000 11.415000 1.600000 ;
      RECT  7.905000 1.600000  8.195000 1.645000 ;
      RECT  8.365000 1.075000  8.655000 1.120000 ;
      RECT  8.365000 1.260000  8.655000 1.305000 ;
      RECT  8.365000 1.755000  8.655000 1.800000 ;
      RECT  8.365000 1.940000  8.655000 1.985000 ;
      RECT 11.125000 1.415000 11.415000 1.460000 ;
      RECT 11.125000 1.600000 11.415000 1.645000 ;
  END
END sky130_fd_sc_hd__sdfbbn_2
MACRO sky130_fd_sc_hd__a222oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a222oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615000 1.000000 2.925000 1.330000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095000 1.000000 3.435000 1.330000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.135000 1.000000 2.445000 1.330000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655000 1.000000 1.965000 1.330000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.000000 0.545000 1.315000 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.715000 1.000000 1.085000 1.315000 ;
    END
  END C2
  PIN Y
    ANTENNADIFFAREA  0.897600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.255000 0.425000 0.645000 ;
        RECT 0.095000 0.645000 2.645000 0.815000 ;
        RECT 0.095000 1.485000 0.425000 1.500000 ;
        RECT 0.095000 1.500000 1.425000 1.670000 ;
        RECT 0.095000 1.670000 0.425000 1.680000 ;
        RECT 0.095000 1.680000 0.345000 2.255000 ;
        RECT 0.095000 2.255000 0.425000 2.465000 ;
        RECT 1.015000 1.670000 1.185000 1.830000 ;
        RECT 1.255000 0.815000 1.480000 1.330000 ;
        RECT 1.255000 1.330000 1.425000 1.500000 ;
        RECT 2.315000 0.295000 2.645000 0.645000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.680000 0.240000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.515000  1.875000 0.845000 2.075000 ;
      RECT 0.595000  2.075000 0.765000 2.295000 ;
      RECT 0.595000  2.295000 2.185000 2.465000 ;
      RECT 0.875000  0.085000 1.605000 0.465000 ;
      RECT 1.515000  1.825000 2.015000 1.965000 ;
      RECT 1.515000  1.965000 1.970000 1.970000 ;
      RECT 1.515000  1.970000 1.935000 1.980000 ;
      RECT 1.515000  1.980000 1.915000 1.995000 ;
      RECT 1.845000  1.655000 3.595000 1.670000 ;
      RECT 1.845000  1.670000 2.685000 1.735000 ;
      RECT 1.845000  1.735000 2.605000 1.825000 ;
      RECT 2.015000  2.135000 2.185000 2.295000 ;
      RECT 2.355000  1.500000 3.595000 1.655000 ;
      RECT 2.355000  1.825000 2.605000 2.255000 ;
      RECT 2.355000  2.255000 2.685000 2.465000 ;
      RECT 2.775000  1.905000 3.105000 2.075000 ;
      RECT 2.855000  2.075000 3.025000 2.635000 ;
      RECT 3.220000  1.670000 3.595000 1.735000 ;
      RECT 3.255000  0.085000 3.585000 0.815000 ;
      RECT 3.255000  2.255000 3.595000 2.465000 ;
      RECT 3.335000  1.735000 3.595000 2.255000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a222oi_1
MACRO sky130_fd_sc_hd__o221ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.430000 1.075000 3.760000 1.445000 ;
        RECT 3.430000 1.445000 4.815000 1.615000 ;
        RECT 4.645000 1.075000 5.435000 1.275000 ;
        RECT 4.645000 1.275000 4.815000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.980000 1.075000 4.475000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 1.075000 2.035000 1.445000 ;
        RECT 1.020000 1.445000 3.260000 1.615000 ;
        RECT 2.930000 1.075000 3.260000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.205000 1.075000 2.760000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.435000 1.275000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.520000 0.645000 0.850000 0.865000 ;
        RECT 0.560000 1.445000 0.850000 1.785000 ;
        RECT 0.560000 1.785000 4.350000 1.955000 ;
        RECT 0.560000 1.955000 0.810000 2.465000 ;
        RECT 0.605000 0.865000 0.850000 1.445000 ;
        RECT 2.340000 1.955000 2.590000 2.125000 ;
        RECT 4.100000 1.955000 4.350000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.100000  0.255000 1.270000 0.475000 ;
      RECT 0.100000  0.475000 0.350000 0.895000 ;
      RECT 0.140000  1.455000 0.390000 2.635000 ;
      RECT 0.980000  2.125000 1.750000 2.635000 ;
      RECT 1.020000  0.475000 1.270000 0.645000 ;
      RECT 1.020000  0.645000 3.050000 0.905000 ;
      RECT 1.460000  0.255000 3.550000 0.475000 ;
      RECT 1.920000  2.125000 2.170000 2.295000 ;
      RECT 1.920000  2.295000 3.010000 2.465000 ;
      RECT 2.760000  2.125000 3.010000 2.295000 ;
      RECT 3.180000  2.125000 3.510000 2.635000 ;
      RECT 3.220000  0.475000 3.550000 0.735000 ;
      RECT 3.220000  0.735000 5.230000 0.905000 ;
      RECT 3.680000  2.125000 3.930000 2.295000 ;
      RECT 3.680000  2.295000 4.770000 2.465000 ;
      RECT 3.720000  0.085000 3.890000 0.555000 ;
      RECT 4.060000  0.255000 4.390000 0.725000 ;
      RECT 4.060000  0.725000 5.230000 0.735000 ;
      RECT 4.520000  1.785000 4.770000 2.295000 ;
      RECT 4.560000  0.085000 4.730000 0.555000 ;
      RECT 4.900000  0.255000 5.230000 0.725000 ;
      RECT 4.985000  1.455000 5.190000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__o221ai_2
MACRO sky130_fd_sc_hd__o221ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675000 1.075000 3.135000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.165000 1.075000 2.505000 1.245000 ;
        RECT 2.295000 1.245000 2.505000 1.445000 ;
        RECT 2.295000 1.445000 2.675000 1.615000 ;
        RECT 2.465000 1.615000 2.675000 2.405000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.995000 1.355000 1.325000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 1.985000 1.325000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.465000 1.325000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.899000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.365000 0.345000 0.645000 ;
        RECT 0.085000 0.645000 0.840000 0.825000 ;
        RECT 0.085000 1.495000 2.125000 1.705000 ;
        RECT 0.085000 1.705000 0.365000 2.465000 ;
        RECT 0.635000 0.825000 0.840000 1.495000 ;
        RECT 1.735000 1.705000 2.125000 1.785000 ;
        RECT 1.735000 1.785000 2.245000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.515000  0.305000 1.775000 0.475000 ;
      RECT 0.550000  1.875000 1.340000 2.635000 ;
      RECT 1.010000  0.645000 2.220000 0.695000 ;
      RECT 1.010000  0.695000 3.135000 0.825000 ;
      RECT 1.945000  0.280000 2.220000 0.645000 ;
      RECT 2.105000  0.825000 3.135000 0.865000 ;
      RECT 2.455000  0.085000 2.625000 0.525000 ;
      RECT 2.795000  0.280000 3.135000 0.695000 ;
      RECT 2.875000  1.455000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o221ai_1
MACRO sky130_fd_sc_hd__o221ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.965000 1.075000 6.295000 1.445000 ;
        RECT 5.965000 1.445000 8.420000 1.615000 ;
        RECT 8.155000 1.075000 9.575000 1.275000 ;
        RECT 8.155000 1.275000 8.420000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.475000 1.075000 7.885000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.360000 1.075000 4.505000 1.275000 ;
        RECT 4.335000 1.275000 4.505000 1.495000 ;
        RECT 4.335000 1.495000 5.795000 1.665000 ;
        RECT 5.465000 1.075000 5.795000 1.495000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675000 0.995000 5.285000 1.325000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.750000 1.275000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.645000 2.125000 0.865000 ;
        RECT 0.575000 1.445000 4.165000 1.615000 ;
        RECT 0.575000 1.615000 0.825000 2.465000 ;
        RECT 1.415000 1.615000 2.125000 1.955000 ;
        RECT 1.415000 1.955000 1.665000 2.465000 ;
        RECT 1.920000 0.865000 2.125000 1.445000 ;
        RECT 3.995000 1.615000 4.165000 1.835000 ;
        RECT 3.995000 1.835000 7.725000 1.955000 ;
        RECT 3.995000 1.955000 6.885000 2.005000 ;
        RECT 3.995000 2.005000 4.285000 2.125000 ;
        RECT 4.875000 2.005000 5.085000 2.125000 ;
        RECT 5.965000 1.785000 7.725000 1.835000 ;
        RECT 6.675000 2.005000 6.885000 2.125000 ;
        RECT 7.475000 1.955000 7.725000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.115000  0.255000 5.585000 0.475000 ;
      RECT 0.115000  0.475000 0.365000 0.895000 ;
      RECT 0.155000  1.485000 0.405000 2.635000 ;
      RECT 0.995000  1.825000 1.245000 2.635000 ;
      RECT 1.835000  2.125000 2.605000 2.635000 ;
      RECT 2.315000  0.645000 6.085000 0.735000 ;
      RECT 2.315000  0.735000 9.445000 0.820000 ;
      RECT 2.775000  1.785000 3.825000 1.955000 ;
      RECT 2.775000  1.955000 3.025000 2.465000 ;
      RECT 3.195000  2.125000 3.445000 2.635000 ;
      RECT 3.615000  1.955000 3.825000 2.295000 ;
      RECT 3.615000  2.295000 5.585000 2.465000 ;
      RECT 4.455000  2.175000 4.705000 2.295000 ;
      RECT 5.255000  2.175000 5.585000 2.295000 ;
      RECT 5.465000  0.820000 9.445000 0.905000 ;
      RECT 5.755000  0.255000 6.085000 0.645000 ;
      RECT 5.755000  2.175000 6.005000 2.635000 ;
      RECT 6.175000  2.175000 6.505000 2.295000 ;
      RECT 6.175000  2.295000 8.145000 2.465000 ;
      RECT 6.255000  0.085000 6.425000 0.555000 ;
      RECT 6.595000  0.255000 6.925000 0.725000 ;
      RECT 6.595000  0.725000 7.765000 0.735000 ;
      RECT 7.055000  2.125000 7.305000 2.295000 ;
      RECT 7.095000  0.085000 7.265000 0.555000 ;
      RECT 7.435000  0.255000 7.765000 0.725000 ;
      RECT 7.895000  1.785000 8.985000 1.955000 ;
      RECT 7.895000  1.955000 8.145000 2.295000 ;
      RECT 7.935000  0.085000 8.105000 0.555000 ;
      RECT 8.275000  0.255000 8.605000 0.725000 ;
      RECT 8.275000  0.725000 9.445000 0.735000 ;
      RECT 8.315000  2.125000 8.565000 2.635000 ;
      RECT 8.735000  1.445000 8.985000 1.785000 ;
      RECT 8.735000  1.955000 8.985000 2.465000 ;
      RECT 8.775000  0.085000 8.945000 0.555000 ;
      RECT 9.115000  0.255000 9.445000 0.725000 ;
      RECT 9.155000  1.445000 9.405000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__o221ai_4
MACRO sky130_fd_sc_hd__fill_8
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.130000 -0.120000 0.350000 0.050000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__fill_8
MACRO sky130_fd_sc_hd__fill_4
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.175000 -0.060000 0.285000 0.060000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__fill_4
MACRO sky130_fd_sc_hd__fill_1
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.055000 0.260000 0.055000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__fill_1
MACRO sky130_fd_sc_hd__fill_2
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.920000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.920000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155000 -0.050000 0.315000 0.060000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.110000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.920000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.920000 0.085000 ;
      RECT 0.000000  2.635000 0.920000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
  END
END sky130_fd_sc_hd__fill_2
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.852000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.400000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.280000 0.280000 2.540000 0.735000 ;
        RECT 2.280000 0.735000 9.025000 0.905000 ;
        RECT 2.315000 1.495000 9.025000 1.720000 ;
        RECT 2.315000 1.720000 7.685000 1.735000 ;
        RECT 2.315000 1.735000 2.540000 2.460000 ;
        RECT 3.140000 0.280000 3.400000 0.735000 ;
        RECT 3.140000 1.735000 3.400000 2.460000 ;
        RECT 4.000000 0.280000 4.260000 0.735000 ;
        RECT 4.000000 1.735000 4.260000 2.460000 ;
        RECT 4.845000 0.280000 5.120000 0.735000 ;
        RECT 4.860000 1.735000 5.120000 2.460000 ;
        RECT 5.705000 0.280000 5.965000 0.735000 ;
        RECT 5.705000 1.735000 5.965000 2.460000 ;
        RECT 6.565000 0.280000 6.825000 0.735000 ;
        RECT 6.565000 1.735000 6.825000 2.460000 ;
        RECT 7.425000 0.280000 7.685000 0.735000 ;
        RECT 7.425000 1.735000 7.685000 2.460000 ;
        RECT 7.860000 0.905000 9.025000 1.495000 ;
        RECT 8.295000 0.280000 8.555000 0.735000 ;
        RECT 8.295000 1.720000 8.585000 2.460000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.495000 0.425000 2.465000 ;
      LAYER mcon ;
        RECT 0.175000 2.125000 0.345000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.955000 1.495000 1.285000 2.465000 ;
      LAYER mcon ;
        RECT 1.035000 2.125000 1.205000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.815000 1.495000 2.145000 2.465000 ;
      LAYER mcon ;
        RECT 1.890000 2.125000 2.060000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.710000 1.905000 2.970000 2.465000 ;
      LAYER mcon ;
        RECT 2.740000 2.125000 2.910000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.570000 1.905000 3.830000 2.465000 ;
      LAYER mcon ;
        RECT 3.620000 2.125000 3.790000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.430000 1.905000 4.690000 2.465000 ;
      LAYER mcon ;
        RECT 4.480000 2.125000 4.650000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.290000 1.905000 5.535000 2.465000 ;
      LAYER mcon ;
        RECT 5.335000 2.125000 5.505000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.150000 1.905000 6.395000 2.465000 ;
      LAYER mcon ;
        RECT 6.195000 2.125000 6.365000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.010000 1.905000 7.255000 2.465000 ;
      LAYER mcon ;
        RECT 7.050000 2.125000 7.220000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.870000 1.905000 8.125000 2.465000 ;
      LAYER mcon ;
        RECT 7.900000 2.125000 8.070000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.755000 1.890000 9.025000 2.465000 ;
      LAYER mcon ;
        RECT 8.780000 2.125000 8.950000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 9.130000 2.340000 ;
        RECT 0.115000 2.080000 0.405000 2.140000 ;
        RECT 0.975000 2.080000 1.265000 2.140000 ;
        RECT 1.830000 2.080000 2.120000 2.140000 ;
        RECT 2.680000 2.080000 2.970000 2.140000 ;
        RECT 3.560000 2.080000 3.850000 2.140000 ;
        RECT 4.420000 2.080000 4.710000 2.140000 ;
        RECT 5.275000 2.080000 5.565000 2.140000 ;
        RECT 6.135000 2.080000 6.425000 2.140000 ;
        RECT 6.990000 2.080000 7.280000 2.140000 ;
        RECT 7.840000 2.080000 8.130000 2.140000 ;
        RECT 8.720000 2.080000 9.010000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.085000  0.085000 0.390000 0.595000 ;
      RECT 0.595000  0.265000 0.820000 1.075000 ;
      RECT 0.595000  1.075000 7.690000 1.325000 ;
      RECT 0.595000  1.325000 0.785000 2.465000 ;
      RECT 0.990000  0.085000 1.250000 0.610000 ;
      RECT 1.430000  0.265000 1.680000 1.075000 ;
      RECT 1.455000  1.325000 1.645000 2.460000 ;
      RECT 1.850000  0.085000 2.110000 0.645000 ;
      RECT 2.710000  0.085000 2.970000 0.565000 ;
      RECT 3.570000  0.085000 3.830000 0.565000 ;
      RECT 4.430000  0.085000 4.675000 0.565000 ;
      RECT 5.290000  0.085000 5.535000 0.565000 ;
      RECT 6.145000  0.085000 6.395000 0.565000 ;
      RECT 7.005000  0.085000 7.255000 0.565000 ;
      RECT 7.865000  0.085000 8.125000 0.565000 ;
      RECT 8.725000  0.085000 9.025000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_16
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.745000 0.785000 1.240000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.383400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 0.255000 1.245000 0.655000 ;
        RECT 1.040000 0.655000 1.725000 0.825000 ;
        RECT 1.060000 1.750000 1.725000 1.970000 ;
        RECT 1.060000 1.970000 1.245000 2.435000 ;
        RECT 1.385000 0.825000 1.725000 1.750000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.855000 0.855000 2.465000 ;
      LAYER mcon ;
        RECT 0.610000 2.125000 0.780000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.415000 2.140000 1.750000 2.465000 ;
      LAYER mcon ;
        RECT 1.495000 2.140000 1.665000 2.310000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 1.770000 2.340000 ;
        RECT 0.550000 2.080000 0.840000 2.140000 ;
        RECT 1.435000 2.080000 1.725000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.410000 ;
      RECT 0.085000  1.410000 1.215000 1.580000 ;
      RECT 0.085000  1.580000 0.355000 2.435000 ;
      RECT 0.555000  0.085000 0.830000 0.565000 ;
      RECT 0.965000  0.995000 1.215000 1.410000 ;
      RECT 1.415000  0.085000 1.750000 0.485000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_2
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.755000 0.775000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.795200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.345000 1.305000 0.735000 ;
        RECT 1.010000 0.735000 2.660000 0.905000 ;
        RECT 1.025000 1.835000 2.165000 1.965000 ;
        RECT 1.025000 1.965000 1.390000 1.970000 ;
        RECT 1.025000 1.970000 1.385000 1.975000 ;
        RECT 1.025000 1.975000 1.370000 1.980000 ;
        RECT 1.025000 1.980000 1.330000 2.000000 ;
        RECT 1.025000 2.000000 1.325000 2.005000 ;
        RECT 1.025000 2.005000 1.265000 2.465000 ;
        RECT 1.185000 1.825000 2.165000 1.835000 ;
        RECT 1.195000 1.820000 2.165000 1.825000 ;
        RECT 1.205000 1.815000 2.165000 1.820000 ;
        RECT 1.215000 1.805000 2.165000 1.815000 ;
        RECT 1.245000 1.785000 2.165000 1.805000 ;
        RECT 1.270000 1.750000 2.165000 1.785000 ;
        RECT 1.905000 0.345000 2.165000 0.735000 ;
        RECT 1.905000 1.415000 2.660000 1.585000 ;
        RECT 1.905000 1.585000 2.165000 1.750000 ;
        RECT 1.935000 1.965000 2.165000 2.465000 ;
        RECT 2.255000 0.905000 2.660000 1.415000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.835000 0.855000 2.465000 ;
      LAYER mcon ;
        RECT 0.610000 2.125000 0.780000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.435000 2.140000 1.765000 2.465000 ;
        RECT 2.335000 1.765000 2.620000 2.465000 ;
      LAYER mcon ;
        RECT 1.495000 2.140000 1.665000 2.310000 ;
        RECT 2.375000 2.125000 2.545000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 2.690000 2.340000 ;
        RECT 0.550000 2.080000 0.840000 2.140000 ;
        RECT 1.435000 2.080000 1.725000 2.140000 ;
        RECT 2.315000 2.080000 2.605000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.255000 0.385000 0.585000 ;
      RECT 0.085000  0.585000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 1.115000 1.665000 ;
      RECT 0.085000  1.665000 0.355000 2.465000 ;
      RECT 0.555000  0.085000 0.830000 0.565000 ;
      RECT 0.945000  1.075000 2.085000 1.245000 ;
      RECT 0.945000  1.245000 1.115000 1.495000 ;
      RECT 1.475000  0.085000 1.730000 0.565000 ;
      RECT 2.335000  0.085000 2.615000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_4
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.426000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 0.400000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.590400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 0.280000 1.680000 0.735000 ;
        RECT 1.420000 0.735000 4.730000 0.905000 ;
        RECT 1.420000 1.495000 4.730000 1.735000 ;
        RECT 1.420000 1.735000 1.680000 2.460000 ;
        RECT 2.280000 0.280000 2.540000 0.735000 ;
        RECT 2.280000 1.735000 2.540000 2.460000 ;
        RECT 3.140000 0.280000 3.400000 0.735000 ;
        RECT 3.140000 1.735000 3.400000 2.460000 ;
        RECT 3.760000 0.905000 4.730000 1.495000 ;
        RECT 4.000000 0.280000 4.260000 0.735000 ;
        RECT 4.000000 1.735000 4.260000 2.460000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.525000 0.390000 2.465000 ;
      LAYER mcon ;
        RECT 0.175000 2.125000 0.345000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.990000 1.525000 1.250000 2.465000 ;
      LAYER mcon ;
        RECT 1.035000 2.125000 1.205000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.850000 1.905000 2.110000 2.465000 ;
      LAYER mcon ;
        RECT 1.890000 2.125000 2.060000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.710000 1.905000 2.970000 2.465000 ;
      LAYER mcon ;
        RECT 2.740000 2.125000 2.910000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.570000 1.905000 3.830000 2.465000 ;
      LAYER mcon ;
        RECT 3.620000 2.125000 3.790000 2.295000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.430000 1.905000 4.725000 2.465000 ;
      LAYER mcon ;
        RECT 4.480000 2.125000 4.650000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 4.990000 2.340000 ;
        RECT 0.115000 2.080000 0.405000 2.140000 ;
        RECT 0.975000 2.080000 1.265000 2.140000 ;
        RECT 1.830000 2.080000 2.120000 2.140000 ;
        RECT 2.680000 2.080000 2.970000 2.140000 ;
        RECT 3.560000 2.080000 3.850000 2.140000 ;
        RECT 4.420000 2.080000 4.710000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.145000  0.085000 0.390000 0.545000 ;
      RECT 0.570000  0.265000 0.820000 1.075000 ;
      RECT 0.570000  1.075000 3.590000 1.325000 ;
      RECT 0.570000  1.325000 0.820000 2.460000 ;
      RECT 0.990000  0.085000 1.250000 0.610000 ;
      RECT 1.850000  0.085000 2.110000 0.565000 ;
      RECT 2.710000  0.085000 2.970000 0.565000 ;
      RECT 3.570000  0.085000 3.830000 0.565000 ;
      RECT 4.430000  0.085000 4.730000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_8
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.196500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.985000 1.275000 1.355000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.345000 0.760000 ;
        RECT 0.085000 0.760000 0.255000 1.560000 ;
        RECT 0.085000 1.560000 0.355000 2.465000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.875000 0.855000 2.465000 ;
      LAYER mcon ;
        RECT 0.610000 2.125000 0.780000 2.295000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 1.310000 2.340000 ;
        RECT 0.550000 2.080000 0.840000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.425000  1.060000 0.710000 1.390000 ;
      RECT 0.525000  0.085000 0.855000 0.465000 ;
      RECT 0.540000  0.635000 1.205000 0.805000 ;
      RECT 0.540000  0.805000 0.710000 1.060000 ;
      RECT 0.540000  1.390000 0.710000 1.535000 ;
      RECT 0.540000  1.535000 1.205000 1.705000 ;
      RECT 1.035000  0.255000 1.205000 0.635000 ;
      RECT 1.035000  1.705000 1.205000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_1
MACRO sky130_fd_sc_hd__a21oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.815000 0.995000 1.425000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.035000 0.645000 1.495000 ;
        RECT 0.145000 1.495000 1.930000 1.675000 ;
        RECT 1.605000 1.075000 1.935000 1.245000 ;
        RECT 1.605000 1.245000 1.930000 1.495000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.800000 0.995000 3.075000 1.625000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.627500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 0.255000 1.300000 0.615000 ;
        RECT 0.955000 0.615000 2.615000 0.785000 ;
        RECT 2.295000 0.255000 2.615000 0.615000 ;
        RECT 2.315000 0.785000 2.615000 2.115000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.100000  0.085000 0.395000 0.865000 ;
      RECT 0.110000  1.855000 2.145000 2.025000 ;
      RECT 0.110000  2.025000 1.220000 2.105000 ;
      RECT 0.110000  2.105000 0.370000 2.465000 ;
      RECT 0.540000  2.275000 0.870000 2.635000 ;
      RECT 1.050000  2.105000 1.220000 2.465000 ;
      RECT 1.475000  2.195000 1.645000 2.635000 ;
      RECT 1.760000  0.085000 2.090000 0.445000 ;
      RECT 1.815000  2.025000 2.145000 2.285000 ;
      RECT 1.815000  2.285000 3.090000 2.465000 ;
      RECT 2.785000  1.795000 3.090000 2.285000 ;
      RECT 2.795000  0.085000 3.125000 0.825000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a21oi_2
MACRO sky130_fd_sc_hd__a21oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.850000 0.995000 1.265000 1.325000 ;
        RECT 1.035000 0.375000 1.265000 0.995000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 0.995000 1.740000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.675000 0.335000 1.325000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.447000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.495000 0.680000 1.685000 ;
        RECT 0.095000 1.685000 0.370000 2.455000 ;
        RECT 0.505000 0.645000 0.835000 0.825000 ;
        RECT 0.505000 0.825000 0.680000 1.495000 ;
        RECT 0.610000 0.265000 0.835000 0.645000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.110000  0.085000 0.440000 0.475000 ;
      RECT 0.540000  1.855000 1.745000 2.025000 ;
      RECT 0.540000  2.025000 0.870000 2.455000 ;
      RECT 0.850000  1.525000 1.745000 1.855000 ;
      RECT 1.040000  2.195000 1.235000 2.635000 ;
      RECT 1.415000  2.025000 1.745000 2.455000 ;
      RECT 1.445000  0.085000 1.745000 0.815000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__a21oi_1
MACRO sky130_fd_sc_hd__a21oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.565000 1.065000 4.000000 1.310000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.050000 1.065000 2.395000 1.480000 ;
        RECT 2.050000 1.480000 5.470000 1.705000 ;
        RECT 4.225000 1.075000 5.470000 1.480000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.400000 1.035000 ;
        RECT 0.090000 1.035000 1.430000 1.415000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.288000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 1.585000 1.880000 1.705000 ;
        RECT 0.580000 1.705000 1.745000 2.035000 ;
        RECT 0.595000 0.370000 0.785000 0.615000 ;
        RECT 0.595000 0.615000 1.645000 0.695000 ;
        RECT 0.595000 0.695000 3.905000 0.865000 ;
        RECT 1.455000 0.255000 1.645000 0.615000 ;
        RECT 1.600000 0.865000 3.905000 0.895000 ;
        RECT 1.600000 0.895000 1.880000 1.585000 ;
        RECT 2.275000 0.675000 3.905000 0.695000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.805000 ;
      RECT 0.180000  1.795000 0.375000 2.215000 ;
      RECT 0.180000  2.215000 2.115000 2.465000 ;
      RECT 0.955000  0.085000 1.285000 0.445000 ;
      RECT 0.955000  2.205000 2.115000 2.215000 ;
      RECT 1.835000  0.085000 2.115000 0.525000 ;
      RECT 1.915000  1.875000 5.625000 2.105000 ;
      RECT 1.915000  2.105000 2.115000 2.205000 ;
      RECT 2.285000  0.255000 4.335000 0.505000 ;
      RECT 2.285000  2.275000 2.615000 2.635000 ;
      RECT 2.785000  2.105000 2.975000 2.465000 ;
      RECT 3.145000  2.275000 3.475000 2.635000 ;
      RECT 3.645000  2.105000 3.835000 2.465000 ;
      RECT 4.005000  2.275000 4.335000 2.635000 ;
      RECT 4.075000  0.505000 4.335000 0.735000 ;
      RECT 4.075000  0.735000 5.195000 0.905000 ;
      RECT 4.505000  0.085000 4.695000 0.565000 ;
      RECT 4.505000  2.105000 4.685000 2.465000 ;
      RECT 4.865000  0.255000 5.195000 0.735000 ;
      RECT 4.865000  2.275000 5.195000 2.635000 ;
      RECT 5.365000  0.085000 5.625000 0.885000 ;
      RECT 5.365000  2.105000 5.625000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__a21oi_4
MACRO sky130_fd_sc_hd__o31a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.140000 1.055000 5.470000 1.360000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.265000 1.055000 4.970000 1.360000 ;
        RECT 4.680000 1.360000 4.970000 1.530000 ;
        RECT 4.680000 1.530000 6.355000 1.700000 ;
        RECT 5.640000 1.055000 6.355000 1.530000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 1.055000 4.095000 1.360000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.780000 1.055000 3.575000 1.355000 ;
        RECT 2.780000 1.355000 3.150000 1.695000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.715000 1.765000 0.885000 ;
        RECT 0.085000 0.885000 0.735000 1.460000 ;
        RECT 0.085000 1.460000 1.750000 1.665000 ;
        RECT 0.680000 0.255000 0.895000 0.655000 ;
        RECT 0.680000 0.655000 1.765000 0.715000 ;
        RECT 0.680000 1.665000 0.895000 2.465000 ;
        RECT 1.565000 0.255000 1.765000 0.655000 ;
        RECT 1.565000 1.665000 1.750000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125000 -0.085000 0.295000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  0.085000 0.510000 0.545000 ;
      RECT 0.085000  1.835000 0.510000 2.635000 ;
      RECT 0.905000  1.055000 2.610000 1.290000 ;
      RECT 1.065000  0.085000 1.395000 0.485000 ;
      RECT 1.065000  1.835000 1.395000 2.635000 ;
      RECT 1.920000  1.460000 2.250000 2.635000 ;
      RECT 1.935000  0.085000 2.250000 0.885000 ;
      RECT 2.440000  0.255000 3.570000 0.465000 ;
      RECT 2.440000  0.635000 3.210000 0.885000 ;
      RECT 2.440000  0.885000 2.610000 1.055000 ;
      RECT 2.440000  1.290000 2.610000 1.870000 ;
      RECT 2.440000  1.870000 4.090000 2.070000 ;
      RECT 2.440000  2.070000 2.610000 2.465000 ;
      RECT 2.780000  2.240000 3.110000 2.635000 ;
      RECT 3.320000  1.530000 4.510000 1.700000 ;
      RECT 3.380000  0.465000 3.570000 0.635000 ;
      RECT 3.380000  0.635000 6.355000 0.885000 ;
      RECT 3.760000  0.085000 4.090000 0.445000 ;
      RECT 3.760000  2.070000 4.090000 2.465000 ;
      RECT 4.260000  0.255000 4.430000 0.635000 ;
      RECT 4.260000  1.700000 4.510000 2.465000 ;
      RECT 4.600000  0.085000 4.930000 0.445000 ;
      RECT 4.680000  1.870000 5.720000 2.070000 ;
      RECT 4.680000  2.070000 4.850000 2.465000 ;
      RECT 5.020000  2.240000 5.350000 2.635000 ;
      RECT 5.100000  0.255000 5.270000 0.635000 ;
      RECT 5.440000  0.085000 5.770000 0.445000 ;
      RECT 5.520000  2.070000 5.720000 2.465000 ;
      RECT 5.890000  1.870000 6.355000 2.465000 ;
      RECT 5.940000  0.255000 6.355000 0.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.125000 4.455000 2.295000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.125000 6.295000 2.295000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 4.225000 2.095000 4.515000 2.140000 ;
      RECT 4.225000 2.140000 6.355000 2.280000 ;
      RECT 4.225000 2.280000 4.515000 2.325000 ;
      RECT 6.065000 2.095000 6.355000 2.140000 ;
      RECT 6.065000 2.280000 6.355000 2.325000 ;
  END
END sky130_fd_sc_hd__o31a_4
MACRO sky130_fd_sc_hd__o31a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.905000 0.995000 1.295000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 0.995000 1.725000 1.325000 ;
        RECT 1.525000 1.325000 1.725000 2.125000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 0.995000 2.175000 2.125000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.390000 0.995000 2.795000 1.325000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.594000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.265000 0.525000 0.825000 ;
        RECT 0.085000 0.825000 0.395000 1.835000 ;
        RECT 0.085000 1.835000 0.525000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.565000  0.995000 0.735000 1.445000 ;
      RECT 0.565000  1.445000 1.355000 1.615000 ;
      RECT 0.695000  0.085000 1.145000 0.825000 ;
      RECT 0.700000  1.785000 1.015000 2.635000 ;
      RECT 1.185000  1.615000 1.355000 2.295000 ;
      RECT 1.185000  2.295000 2.615000 2.465000 ;
      RECT 1.315000  0.255000 1.485000 0.655000 ;
      RECT 1.315000  0.655000 2.475000 0.825000 ;
      RECT 1.655000  0.085000 2.075000 0.485000 ;
      RECT 2.245000  0.255000 2.475000 0.655000 ;
      RECT 2.365000  1.495000 3.135000 1.665000 ;
      RECT 2.365000  1.665000 2.615000 2.295000 ;
      RECT 2.645000  0.255000 3.135000 0.825000 ;
      RECT 2.795000  1.835000 3.125000 2.635000 ;
      RECT 2.965000  0.825000 3.135000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o31a_1
MACRO sky130_fd_sc_hd__o31a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.370000 0.995000 1.760000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 0.995000 2.190000 1.325000 ;
        RECT 1.990000 1.325000 2.190000 2.125000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.390000 0.995000 2.640000 2.125000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855000 0.995000 3.255000 1.325000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.577500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.860000 1.295000 ;
        RECT 0.550000 0.265000 0.990000 0.825000 ;
        RECT 0.550000 0.825000 0.860000 1.075000 ;
        RECT 0.550000 1.295000 0.860000 1.835000 ;
        RECT 0.550000 1.835000 0.990000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 0.380000 0.905000 ;
      RECT 0.085000  1.465000 0.380000 2.635000 ;
      RECT 1.030000  0.995000 1.200000 1.445000 ;
      RECT 1.030000  1.445000 1.820000 1.615000 ;
      RECT 1.160000  0.085000 1.610000 0.825000 ;
      RECT 1.165000  1.785000 1.480000 2.635000 ;
      RECT 1.650000  1.615000 1.820000 2.295000 ;
      RECT 1.650000  2.295000 3.080000 2.465000 ;
      RECT 1.780000  0.255000 1.950000 0.655000 ;
      RECT 1.780000  0.655000 2.940000 0.825000 ;
      RECT 2.120000  0.085000 2.540000 0.485000 ;
      RECT 2.710000  0.255000 2.940000 0.655000 ;
      RECT 2.830000  1.495000 3.595000 1.665000 ;
      RECT 2.830000  1.665000 3.080000 2.295000 ;
      RECT 3.110000  0.255000 3.595000 0.825000 ;
      RECT 3.255000  1.835000 3.590000 2.635000 ;
      RECT 3.425000  0.825000 3.595000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__o31a_2
MACRO sky130_fd_sc_hd__tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tap_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.265000 0.375000 0.810000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.315000 0.845000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.470000 0.375000 2.455000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__tap_1
MACRO sky130_fd_sc_hd__tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tap_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.920000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.920000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.265000 0.835000 0.810000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.775000 0.845000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.470000 0.835000 2.455000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 1.110000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.920000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.920000 0.085000 ;
      RECT 0.000000  2.635000 0.920000 2.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
  END
END sky130_fd_sc_hd__tap_2
MACRO sky130_fd_sc_hd__nand2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 1.075000 1.765000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.845000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.495000 2.215000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 0.655000 2.215000 0.905000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 1.935000 0.905000 2.215000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.255000 0.425000 0.715000 ;
      RECT 0.085000  0.715000 1.185000 0.885000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 0.935000  0.255000 2.105000 0.465000 ;
      RECT 0.935000  0.465000 1.185000 0.715000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.775000  0.465000 2.105000 0.485000 ;
      RECT 1.855000  1.835000 2.110000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2_2
MACRO sky130_fd_sc_hd__nand2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615000 1.075000 4.055000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 1.730000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.495000 3.365000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 1.910000 1.075000 2.445000 1.495000 ;
        RECT 2.195000 0.635000 3.365000 0.805000 ;
        RECT 2.195000 0.805000 2.445000 1.075000 ;
        RECT 2.195000 1.665000 2.525000 2.465000 ;
        RECT 3.035000 1.665000 3.365000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.715000 ;
      RECT 0.090000  0.715000 2.025000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.545000 ;
      RECT 0.935000  0.255000 1.265000 0.715000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.435000  0.085000 1.605000 0.545000 ;
      RECT 1.775000  0.255000 3.785000 0.465000 ;
      RECT 1.775000  0.465000 2.025000 0.715000 ;
      RECT 1.855000  1.835000 2.025000 2.635000 ;
      RECT 2.695000  1.835000 2.865000 2.635000 ;
      RECT 3.535000  0.465000 3.785000 0.885000 ;
      RECT 3.535000  1.835000 3.785000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2_4
MACRO sky130_fd_sc_hd__nand2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.290000 1.075000 6.305000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.510000 1.075000 3.365000 1.295000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.862000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.465000 6.725000 1.665000 ;
        RECT 0.515000 1.665000 0.845000 2.465000 ;
        RECT 1.355000 1.665000 1.685000 2.465000 ;
        RECT 2.195000 1.665000 2.525000 2.465000 ;
        RECT 3.035000 1.665000 3.365000 2.465000 ;
        RECT 3.640000 1.075000 4.120000 1.465000 ;
        RECT 3.875000 0.655000 6.725000 0.905000 ;
        RECT 3.875000 0.905000 4.120000 1.075000 ;
        RECT 3.875000 1.665000 4.205000 2.465000 ;
        RECT 4.715000 1.665000 5.045000 2.465000 ;
        RECT 5.555000 1.665000 5.885000 2.465000 ;
        RECT 6.395000 1.665000 6.725000 2.465000 ;
        RECT 6.475000 0.905000 6.725000 1.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.735000 ;
      RECT 0.090000  0.735000 3.705000 0.905000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 0.595000  0.085000 0.765000 0.565000 ;
      RECT 0.935000  0.255000 1.265000 0.735000 ;
      RECT 1.015000  1.835000 1.185000 2.635000 ;
      RECT 1.435000  0.085000 1.605000 0.565000 ;
      RECT 1.775000  0.255000 2.105000 0.735000 ;
      RECT 1.855000  1.835000 2.025000 2.635000 ;
      RECT 2.275000  0.085000 2.445000 0.565000 ;
      RECT 2.615000  0.255000 2.945000 0.735000 ;
      RECT 2.695000  1.835000 2.865000 2.635000 ;
      RECT 3.115000  0.085000 3.285000 0.565000 ;
      RECT 3.455000  0.255000 7.270000 0.485000 ;
      RECT 3.455000  0.485000 3.705000 0.735000 ;
      RECT 3.535000  1.835000 3.705000 2.635000 ;
      RECT 4.375000  1.835000 4.545000 2.635000 ;
      RECT 5.215000  1.835000 5.385000 2.635000 ;
      RECT 6.055000  1.835000 6.225000 2.635000 ;
      RECT 6.895000  0.485000 7.270000 0.905000 ;
      RECT 6.915000  1.495000 7.270000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2_8
MACRO sky130_fd_sc_hd__nand2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.940000 1.075000 1.275000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.055000 0.430000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 1.485000 0.865000 2.465000 ;
        RECT 0.600000 0.255000 1.295000 0.885000 ;
        RECT 0.600000 0.885000 0.770000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.085000  0.085000 0.395000 0.885000 ;
      RECT 0.085000  1.495000 0.365000 2.635000 ;
      RECT 1.035000  1.495000 1.295000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2_1
MACRO sky130_fd_sc_hd__and4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.325000 2.075000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885000 0.360000 1.235000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 0.355000 1.715000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 0.355000 2.175000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.795000 0.295000 3.135000 0.805000 ;
        RECT 2.795000 2.205000 3.135000 2.465000 ;
        RECT 2.875000 0.805000 3.135000 2.205000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  2.255000 0.425000 2.635000 ;
      RECT 0.170000  0.255000 0.665000 0.585000 ;
      RECT 0.495000  0.585000 0.665000 1.495000 ;
      RECT 0.495000  1.495000 2.685000 1.665000 ;
      RECT 0.595000  1.665000 0.845000 2.465000 ;
      RECT 1.065000  1.915000 1.395000 2.635000 ;
      RECT 1.580000  1.665000 1.830000 2.465000 ;
      RECT 2.295000  1.835000 2.625000 2.635000 ;
      RECT 2.355000  0.085000 2.625000 0.885000 ;
      RECT 2.370000  1.075000 2.700000 1.325000 ;
      RECT 2.370000  1.325000 2.685000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__and4_1
MACRO sky130_fd_sc_hd__and4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.755000 0.330000 2.075000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.890000 0.420000 1.245000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 0.415000 1.720000 1.305000 ;
        RECT 1.420000 1.305000 1.590000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.900000 0.415000 2.160000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.544500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 0.295000 3.065000 0.340000 ;
        RECT 2.735000 0.340000 3.070000 0.805000 ;
        RECT 2.735000 1.495000 3.070000 2.465000 ;
        RECT 2.895000 0.805000 3.070000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  2.255000 0.425000 2.635000 ;
      RECT 0.175000  0.255000 0.670000 0.585000 ;
      RECT 0.500000  0.585000 0.670000 1.495000 ;
      RECT 0.500000  1.495000 2.555000 1.665000 ;
      RECT 0.600000  1.665000 0.850000 2.465000 ;
      RECT 1.070000  1.915000 1.400000 2.635000 ;
      RECT 1.585000  1.665000 1.835000 2.465000 ;
      RECT 2.235000  1.835000 2.565000 2.635000 ;
      RECT 2.330000  0.085000 2.565000 0.890000 ;
      RECT 2.330000  1.075000 2.725000 1.315000 ;
      RECT 2.330000  1.315000 2.555000 1.495000 ;
      RECT 3.245000  1.835000 3.575000 2.635000 ;
      RECT 3.255000  0.085000 3.585000 0.810000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__and4_2
MACRO sky130_fd_sc_hd__and4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.765000 0.330000 1.655000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.840000 0.995000 1.245000 1.325000 ;
        RECT 0.890000 0.420000 1.245000 0.995000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 0.425000 1.700000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.905000 0.730000 2.155000 0.935000 ;
        RECT 1.905000 0.935000 2.075000 1.325000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.535000 0.255000 2.705000 0.640000 ;
        RECT 2.535000 0.640000 4.050000 0.810000 ;
        RECT 2.535000 1.795000 2.785000 2.465000 ;
        RECT 2.615000 1.485000 4.050000 1.655000 ;
        RECT 2.615000 1.655000 2.785000 1.795000 ;
        RECT 3.375000 0.255000 3.545000 0.640000 ;
        RECT 3.375000 1.655000 4.050000 1.745000 ;
        RECT 3.375000 1.745000 3.545000 2.465000 ;
        RECT 3.800000 0.810000 4.050000 1.485000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.105000  1.835000 0.385000 2.635000 ;
      RECT 0.175000  0.255000 0.670000 0.585000 ;
      RECT 0.500000  0.585000 0.670000 1.495000 ;
      RECT 0.500000  1.495000 2.415000 1.665000 ;
      RECT 0.555000  1.665000 0.765000 2.465000 ;
      RECT 0.955000  1.935000 1.285000 2.635000 ;
      RECT 1.455000  1.665000 1.645000 2.465000 ;
      RECT 2.025000  0.085000 2.335000 0.550000 ;
      RECT 2.025000  1.855000 2.355000 2.635000 ;
      RECT 2.245000  1.105000 3.585000 1.305000 ;
      RECT 2.245000  1.305000 2.415000 1.495000 ;
      RECT 2.575000  1.075000 3.585000 1.105000 ;
      RECT 2.875000  0.085000 3.205000 0.470000 ;
      RECT 2.955000  1.835000 3.205000 2.635000 ;
      RECT 3.715000  0.085000 4.045000 0.470000 ;
      RECT 3.715000  1.915000 4.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__and4_4
MACRO sky130_fd_sc_hd__lpflow_bleeder_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_bleeder_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN SHORT
    ANTENNAGATEAREA  0.270000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.275000 1.040000 1.975000 1.730000 ;
    END
  END SHORT
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.285000  0.085000 0.615000 0.870000 ;
      RECT 2.145000  0.540000 2.475000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_bleeder_1
MACRO sky130_fd_sc_hd__a22oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.275000 1.075000 5.685000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.910000 1.075000 7.735000 1.285000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615000 1.075000 4.040000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.895000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 1.445000 3.325000 1.625000 ;
        RECT 0.595000 1.625000 0.805000 2.125000 ;
        RECT 1.395000 1.625000 1.645000 2.125000 ;
        RECT 2.195000 0.645000 5.565000 0.885000 ;
        RECT 2.195000 0.885000 2.445000 1.445000 ;
        RECT 2.235000 1.625000 2.485000 2.125000 ;
        RECT 3.075000 1.625000 3.325000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.090000  1.455000 0.425000 2.295000 ;
      RECT 0.090000  2.295000 4.265000 2.465000 ;
      RECT 0.095000  0.255000 0.425000 0.725000 ;
      RECT 0.095000  0.725000 2.025000 0.905000 ;
      RECT 0.595000  0.085000 0.765000 0.555000 ;
      RECT 0.935000  0.255000 1.265000 0.725000 ;
      RECT 0.975000  1.795000 1.225000 2.295000 ;
      RECT 1.435000  0.085000 1.605000 0.555000 ;
      RECT 1.775000  0.255000 3.785000 0.475000 ;
      RECT 1.775000  0.475000 2.025000 0.725000 ;
      RECT 1.815000  1.795000 2.065000 2.295000 ;
      RECT 2.655000  1.795000 2.905000 2.295000 ;
      RECT 3.495000  1.455000 7.625000 1.625000 ;
      RECT 3.495000  1.625000 4.265000 2.295000 ;
      RECT 3.975000  0.255000 5.985000 0.475000 ;
      RECT 4.435000  1.795000 4.685000 2.635000 ;
      RECT 4.855000  1.625000 5.105000 2.465000 ;
      RECT 5.275000  1.795000 5.525000 2.635000 ;
      RECT 5.695000  1.625000 5.945000 2.465000 ;
      RECT 5.735000  0.475000 5.985000 0.725000 ;
      RECT 5.735000  0.725000 7.665000 0.905000 ;
      RECT 6.115000  1.795000 6.365000 2.635000 ;
      RECT 6.155000  0.085000 6.325000 0.555000 ;
      RECT 6.495000  0.255000 6.825000 0.725000 ;
      RECT 6.535000  1.625000 6.785000 2.465000 ;
      RECT 6.955000  1.795000 7.205000 2.635000 ;
      RECT 6.995000  0.085000 7.165000 0.555000 ;
      RECT 7.335000  0.255000 7.665000 0.725000 ;
      RECT 7.375000  1.625000 7.625000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__a22oi_4
MACRO sky130_fd_sc_hd__a22oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.075000 3.100000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.390000 1.075000 4.500000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.075000 1.700000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 1.075000 0.780000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.141000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.485000 2.160000 1.655000 ;
        RECT 0.095000 1.655000 0.345000 2.465000 ;
        RECT 0.935000 1.655000 1.265000 2.125000 ;
        RECT 1.355000 0.675000 3.045000 0.845000 ;
        RECT 1.775000 1.655000 2.160000 2.125000 ;
        RECT 1.870000 0.845000 2.160000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.095000  0.255000 0.345000 0.680000 ;
      RECT 0.095000  0.680000 1.185000 0.850000 ;
      RECT 0.515000  0.085000 0.845000 0.510000 ;
      RECT 0.515000  1.825000 0.765000 2.295000 ;
      RECT 0.515000  2.295000 2.625000 2.465000 ;
      RECT 1.015000  0.255000 2.105000 0.505000 ;
      RECT 1.015000  0.505000 1.185000 0.680000 ;
      RECT 1.435000  1.825000 1.605000 2.295000 ;
      RECT 2.295000  0.255000 3.385000 0.505000 ;
      RECT 2.375000  1.485000 4.305000 1.655000 ;
      RECT 2.375000  1.655000 2.625000 2.295000 ;
      RECT 2.795000  1.825000 2.965000 2.635000 ;
      RECT 3.135000  1.655000 3.465000 2.465000 ;
      RECT 3.215000  0.505000 3.385000 0.680000 ;
      RECT 3.215000  0.680000 4.375000 0.850000 ;
      RECT 3.555000  0.085000 3.885000 0.510000 ;
      RECT 3.635000  1.825000 3.805000 2.635000 ;
      RECT 3.975000  1.655000 4.305000 2.465000 ;
      RECT 4.055000  0.255000 4.375000 0.680000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__a22oi_2
MACRO sky130_fd_sc_hd__a22oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.490000 0.675000 1.700000 1.075000 ;
        RECT 1.490000 1.075000 1.840000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.010000 0.995000 2.335000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765000 1.075000 1.240000 1.275000 ;
        RECT 0.990000 0.675000 1.240000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.765000 0.575000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.858000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.445000 1.840000 1.495000 ;
        RECT 0.095000 1.495000 2.675000 1.625000 ;
        RECT 0.095000 1.625000 0.425000 2.295000 ;
        RECT 0.095000 2.295000 1.265000 2.465000 ;
        RECT 0.820000 0.255000 2.125000 0.505000 ;
        RECT 0.935000 2.255000 1.265000 2.295000 ;
        RECT 1.615000 1.625000 2.675000 1.665000 ;
        RECT 1.945000 0.505000 2.125000 0.655000 ;
        RECT 1.945000 0.655000 2.675000 0.825000 ;
        RECT 2.505000 0.825000 2.675000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  0.085000 0.545000 0.595000 ;
      RECT 0.595000  1.795000 1.475000 1.835000 ;
      RECT 0.595000  1.835000 2.125000 2.035000 ;
      RECT 0.595000  2.035000 1.210000 2.085000 ;
      RECT 0.595000  2.085000 0.825000 2.125000 ;
      RECT 1.435000  2.255000 1.810000 2.635000 ;
      RECT 1.955000  2.035000 2.125000 2.165000 ;
      RECT 2.305000  0.085000 2.635000 0.485000 ;
      RECT 2.360000  1.855000 2.625000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__a22oi_1
MACRO sky130_fd_sc_hd__nand3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.075000 0.780000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.270000 1.075000 4.480000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.790000 1.075000 6.500000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.635000 2.965000 0.905000 ;
        RECT 1.455000 1.445000 6.505000 1.665000 ;
        RECT 1.455000 1.665000 1.785000 2.465000 ;
        RECT 2.295000 1.665000 3.465000 2.005000 ;
        RECT 2.295000 2.005000 2.625000 2.465000 ;
        RECT 2.795000 0.905000 2.965000 1.075000 ;
        RECT 2.795000 1.075000 3.100000 1.445000 ;
        RECT 3.135000 2.005000 3.465000 2.465000 ;
        RECT 3.975000 1.665000 4.305000 2.465000 ;
        RECT 5.335000 1.665000 5.665000 2.465000 ;
        RECT 6.175000 1.665000 6.505000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.085000  0.255000 0.425000 0.715000 ;
      RECT 0.085000  0.715000 1.285000 0.905000 ;
      RECT 0.085000  0.905000 0.260000 1.445000 ;
      RECT 0.085000  1.445000 0.425000 2.465000 ;
      RECT 0.595000  0.085000 0.845000 0.545000 ;
      RECT 0.595000  1.445000 1.285000 2.635000 ;
      RECT 1.005000  0.905000 1.285000 1.075000 ;
      RECT 1.005000  1.075000 2.625000 1.275000 ;
      RECT 1.035000  0.255000 4.725000 0.465000 ;
      RECT 1.955000  1.835000 2.125000 2.635000 ;
      RECT 2.795000  2.175000 2.965000 2.635000 ;
      RECT 3.135000  0.635000 4.725000 0.715000 ;
      RECT 3.135000  0.715000 6.505000 0.905000 ;
      RECT 3.635000  1.835000 3.805000 2.635000 ;
      RECT 4.475000  1.835000 5.165000 2.635000 ;
      RECT 4.915000  0.085000 5.165000 0.545000 ;
      RECT 5.335000  0.255000 5.665000 0.715000 ;
      RECT 5.835000  0.085000 6.005000 0.545000 ;
      RECT 5.835000  1.835000 6.005000 2.635000 ;
      RECT 6.175000  0.255000 6.505000 0.715000 ;
      RECT 6.675000  0.085000 7.005000 0.905000 ;
      RECT 6.675000  1.445000 7.005000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__nand3b_4
MACRO sky130_fd_sc_hd__nand3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.075000 0.780000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.950000 1.075000 3.140000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.075000 1.740000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.785000 4.050000 1.955000 ;
        RECT 1.060000 1.955000 2.230000 2.005000 ;
        RECT 1.060000 2.005000 1.390000 2.465000 ;
        RECT 1.900000 2.005000 2.230000 2.465000 ;
        RECT 3.260000 0.635000 4.050000 0.905000 ;
        RECT 3.260000 1.955000 4.050000 2.005000 ;
        RECT 3.260000 2.005000 3.510000 2.465000 ;
        RECT 3.850000 0.905000 4.050000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.255000 0.410000 0.655000 ;
      RECT 0.090000  0.655000 0.260000 1.445000 ;
      RECT 0.090000  1.445000 3.650000 1.615000 ;
      RECT 0.090000  1.615000 0.260000 2.065000 ;
      RECT 0.090000  2.065000 0.410000 2.465000 ;
      RECT 0.580000  0.085000 0.890000 0.905000 ;
      RECT 0.580000  1.835000 0.890000 2.635000 ;
      RECT 1.060000  0.255000 1.390000 0.715000 ;
      RECT 1.060000  0.715000 2.750000 0.905000 ;
      RECT 1.560000  0.085000 1.810000 0.545000 ;
      RECT 1.560000  2.175000 1.730000 2.635000 ;
      RECT 2.000000  0.255000 4.050000 0.465000 ;
      RECT 2.000000  0.635000 2.750000 0.715000 ;
      RECT 2.400000  2.175000 2.650000 2.635000 ;
      RECT 2.840000  2.175000 3.090000 2.635000 ;
      RECT 2.920000  0.465000 3.090000 0.905000 ;
      RECT 3.320000  1.075000 3.650000 1.445000 ;
      RECT 3.760000  2.175000 4.050000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__nand3b_2
MACRO sky130_fd_sc_hd__nand3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.425000 0.995000 1.755000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 0.995000 1.235000 1.325000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.732000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.130000 1.495000 2.675000 1.665000 ;
        RECT 1.130000 1.665000 1.460000 2.465000 ;
        RECT 2.085000 0.255000 2.675000 0.485000 ;
        RECT 2.085000 1.665000 2.675000 2.465000 ;
        RECT 2.385000 0.485000 2.675000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.445000 0.510000 0.655000 ;
      RECT 0.085000  0.655000 2.215000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.595000 ;
      RECT 0.085000  1.595000 0.510000 1.925000 ;
      RECT 0.710000  0.085000 1.040000 0.485000 ;
      RECT 0.710000  1.495000 0.960000 2.635000 ;
      RECT 1.630000  1.835000 1.915000 2.635000 ;
      RECT 2.045000  0.825000 2.215000 1.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__nand3b_1
MACRO sky130_fd_sc_hd__nor2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.075000 1.800000 1.275000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.075000 4.975000 1.320000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 3.385000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 2.295000 0.905000 2.625000 1.445000 ;
        RECT 2.295000 1.445000 3.305000 1.745000 ;
        RECT 2.295000 1.745000 2.465000 2.125000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 3.135000 1.745000 3.305000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.905000 ;
      RECT 0.085000  1.455000 2.125000 1.665000 ;
      RECT 0.085000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.865000 2.635000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.035000  1.665000 1.205000 2.465000 ;
      RECT 1.375000  1.835000 1.625000 2.635000 ;
      RECT 1.795000  1.665000 2.125000 2.295000 ;
      RECT 1.795000  2.295000 3.855000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.635000  1.935000 2.965000 2.295000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 2.795000  1.075000 4.275000 1.275000 ;
      RECT 3.475000  1.575000 3.855000 2.295000 ;
      RECT 3.555000  0.085000 3.845000 0.905000 ;
      RECT 4.025000  0.255000 4.355000 0.815000 ;
      RECT 4.025000  0.815000 4.275000 1.075000 ;
      RECT 4.025000  1.275000 4.275000 1.575000 ;
      RECT 4.025000  1.575000 4.355000 2.465000 ;
      RECT 4.525000  0.085000 4.815000 0.905000 ;
      RECT 4.525000  1.495000 4.930000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2b_4
MACRO sky130_fd_sc_hd__nor2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.480000 1.065000 0.920000 1.275000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.600000 1.065000 3.125000 1.275000 ;
        RECT 2.910000 1.275000 3.125000 1.965000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 1.705000 0.895000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 1.415000 0.895000 1.665000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.895000 ;
      RECT 0.085000  1.445000 1.245000 1.655000 ;
      RECT 0.085000  1.655000 0.405000 2.465000 ;
      RECT 0.575000  1.825000 0.825000 2.635000 ;
      RECT 0.995000  1.655000 1.245000 2.295000 ;
      RECT 0.995000  2.295000 2.125000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.835000  1.445000 2.090000 1.890000 ;
      RECT 1.835000  1.890000 2.125000 2.295000 ;
      RECT 1.875000  0.085000 2.045000 0.895000 ;
      RECT 1.875000  1.075000 2.430000 1.245000 ;
      RECT 2.215000  0.725000 2.565000 0.895000 ;
      RECT 2.215000  0.895000 2.430000 1.075000 ;
      RECT 2.260000  1.245000 2.430000 1.445000 ;
      RECT 2.260000  1.445000 2.565000 1.615000 ;
      RECT 2.395000  0.445000 2.565000 0.725000 ;
      RECT 2.395000  1.615000 2.565000 2.460000 ;
      RECT 2.775000  0.085000 3.030000 0.845000 ;
      RECT 2.775000  2.145000 3.025000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2b_2
MACRO sky130_fd_sc_hd__nor2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 1.065000 1.325000 1.325000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.725000 0.325000 1.325000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.235000 0.255000 1.565000 0.725000 ;
        RECT 1.235000 0.725000 2.215000 0.895000 ;
        RECT 1.655000 1.850000 2.215000 2.465000 ;
        RECT 2.035000 0.895000 2.215000 1.850000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.330000  0.370000 0.675000 0.545000 ;
      RECT 0.415000  1.510000 1.705000 1.680000 ;
      RECT 0.415000  1.680000 0.675000 1.905000 ;
      RECT 0.495000  0.545000 0.675000 1.510000 ;
      RECT 0.855000  0.085000 1.065000 0.895000 ;
      RECT 0.875000  1.855000 1.205000 2.635000 ;
      RECT 1.535000  1.075000 1.865000 1.245000 ;
      RECT 1.535000  1.245000 1.705000 1.510000 ;
      RECT 1.735000  0.085000 2.120000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2b_1
MACRO sky130_fd_sc_hd__einvp_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.420000 1.020000 8.195000 1.275000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  1.027500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.330000 1.615000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.870000 0.635000 8.195000 0.850000 ;
        RECT 4.870000 0.850000 5.250000 1.445000 ;
        RECT 4.870000 1.445000 7.720000 1.615000 ;
        RECT 4.870000 1.615000 5.200000 2.125000 ;
        RECT 5.710000 1.615000 6.040000 2.125000 ;
        RECT 6.550000 1.615000 6.880000 2.125000 ;
        RECT 7.390000 1.615000 7.720000 2.125000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.695000 0.825000 ;
      RECT 0.085000  1.785000 0.875000 1.955000 ;
      RECT 0.085000  1.955000 0.345000 2.465000 ;
      RECT 0.500000  0.825000 0.695000 0.995000 ;
      RECT 0.500000  0.995000 4.700000 1.325000 ;
      RECT 0.500000  1.325000 0.875000 1.785000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  2.125000 0.875000 2.635000 ;
      RECT 1.035000  0.255000 1.205000 0.655000 ;
      RECT 1.035000  0.655000 4.700000 0.825000 ;
      RECT 1.075000  1.555000 4.700000 1.725000 ;
      RECT 1.075000  1.725000 1.285000 2.465000 ;
      RECT 1.375000  0.085000 1.705000 0.485000 ;
      RECT 1.455000  1.895000 1.785000 2.635000 ;
      RECT 1.875000  0.255000 2.045000 0.655000 ;
      RECT 1.955000  1.725000 2.125000 2.465000 ;
      RECT 2.215000  0.085000 2.545000 0.485000 ;
      RECT 2.295000  1.895000 2.625000 2.635000 ;
      RECT 2.715000  0.255000 2.885000 0.655000 ;
      RECT 2.795000  1.725000 2.965000 2.465000 ;
      RECT 3.055000  0.085000 3.385000 0.485000 ;
      RECT 3.135000  1.895000 3.465000 2.635000 ;
      RECT 3.555000  0.255000 3.725000 0.655000 ;
      RECT 3.635000  1.725000 3.805000 2.465000 ;
      RECT 3.895000  0.085000 4.235000 0.485000 ;
      RECT 3.975000  1.895000 4.305000 2.635000 ;
      RECT 4.405000  0.255000 8.195000 0.465000 ;
      RECT 4.405000  0.465000 4.700000 0.655000 ;
      RECT 4.475000  1.725000 4.700000 2.295000 ;
      RECT 4.475000  2.295000 8.195000 2.465000 ;
      RECT 5.370000  1.785000 5.540000 2.295000 ;
      RECT 6.210000  1.785000 6.380000 2.295000 ;
      RECT 7.050000  1.785000 7.220000 2.295000 ;
      RECT 7.890000  1.445000 8.195000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
END sky130_fd_sc_hd__einvp_8
MACRO sky130_fd_sc_hd__einvp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.740000 1.020000 4.975000 1.275000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.637500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.330000 1.615000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.190000 0.635000 4.975000 0.850000 ;
        RECT 3.190000 0.850000 3.570000 1.445000 ;
        RECT 3.190000 1.445000 4.360000 1.615000 ;
        RECT 3.190000 1.615000 3.520000 2.125000 ;
        RECT 4.030000 1.615000 4.360000 2.125000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.695000 0.825000 ;
      RECT 0.085000  1.785000 0.875000 1.955000 ;
      RECT 0.085000  1.955000 0.345000 2.465000 ;
      RECT 0.500000  0.825000 0.695000 0.995000 ;
      RECT 0.500000  0.995000 3.020000 1.325000 ;
      RECT 0.500000  1.325000 0.875000 1.785000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  2.125000 0.875000 2.635000 ;
      RECT 1.035000  0.255000 1.205000 0.655000 ;
      RECT 1.035000  0.655000 3.020000 0.825000 ;
      RECT 1.075000  1.555000 2.995000 1.725000 ;
      RECT 1.075000  1.725000 1.285000 2.465000 ;
      RECT 1.375000  0.085000 1.705000 0.485000 ;
      RECT 1.455000  1.895000 1.785000 2.635000 ;
      RECT 1.875000  0.255000 2.045000 0.655000 ;
      RECT 1.955000  1.725000 2.125000 2.465000 ;
      RECT 2.215000  0.085000 2.555000 0.485000 ;
      RECT 2.295000  1.895000 2.655000 2.635000 ;
      RECT 2.735000  0.255000 4.975000 0.465000 ;
      RECT 2.735000  0.465000 3.020000 0.655000 ;
      RECT 2.825000  1.725000 2.995000 2.295000 ;
      RECT 2.825000  2.295000 4.975000 2.465000 ;
      RECT 3.690000  1.785000 3.860000 2.295000 ;
      RECT 4.530000  1.445000 4.975000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__einvp_4
MACRO sky130_fd_sc_hd__einvp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.850000 0.765000 3.135000 1.615000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.354000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.330000 1.615000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.350000 0.595000 2.680000 2.125000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.875000 0.825000 ;
      RECT 0.085000  1.785000 0.875000 1.955000 ;
      RECT 0.085000  1.955000 0.345000 2.465000 ;
      RECT 0.500000  0.825000 0.875000 0.995000 ;
      RECT 0.500000  0.995000 2.180000 1.325000 ;
      RECT 0.500000  1.325000 0.875000 1.785000 ;
      RECT 0.515000  0.085000 0.875000 0.485000 ;
      RECT 0.515000  2.125000 0.875000 2.635000 ;
      RECT 1.045000  0.255000 1.240000 0.655000 ;
      RECT 1.045000  0.655000 2.180000 0.825000 ;
      RECT 1.045000  1.555000 2.155000 1.725000 ;
      RECT 1.045000  1.725000 1.285000 2.465000 ;
      RECT 1.410000  0.085000 1.770000 0.485000 ;
      RECT 1.455000  1.895000 1.785000 2.635000 ;
      RECT 1.940000  0.255000 3.135000 0.425000 ;
      RECT 1.940000  0.425000 2.180000 0.655000 ;
      RECT 1.985000  1.725000 2.155000 2.295000 ;
      RECT 1.985000  2.295000 3.135000 2.465000 ;
      RECT 2.850000  0.425000 3.135000 0.595000 ;
      RECT 2.850000  1.785000 3.135000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__einvp_2
MACRO sky130_fd_sc_hd__einvp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 0.975000 2.215000 1.955000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.223500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.545000 1.725000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.620000 0.255000 2.215000 0.805000 ;
        RECT 1.620000 0.805000 1.795000 2.125000 ;
        RECT 1.620000 2.125000 2.215000 2.465000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 1.450000 0.825000 ;
      RECT 0.085000  1.895000 1.450000 2.065000 ;
      RECT 0.085000  2.065000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 1.450000 0.485000 ;
      RECT 0.515000  2.235000 1.450000 2.635000 ;
      RECT 0.715000  0.825000 1.450000 1.895000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__einvp_1
MACRO sky130_fd_sc_hd__sdfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.460000 1.355000 2.795000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.285000 0.305000  9.615000 0.735000 ;
        RECT  9.285000 0.735000 10.955000 0.905000 ;
        RECT  9.285000 1.505000 10.955000 1.675000 ;
        RECT  9.285000 1.675000  9.615000 2.395000 ;
        RECT 10.135000 0.305000 10.465000 0.735000 ;
        RECT 10.135000 1.675000 10.465000 2.395000 ;
        RECT 10.655000 0.905000 10.955000 1.505000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.535000 1.035000 4.025000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.615000 3.255000 0.785000 ;
        RECT 1.780000 0.785000 1.950000 1.685000 ;
        RECT 2.475000 0.305000 2.650000 0.615000 ;
        RECT 3.085000 0.785000 3.255000 1.115000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.810000 0.805000 ;
      RECT  0.180000  1.795000  0.845000 1.965000 ;
      RECT  0.180000  1.965000  0.350000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.520000  2.135000  0.850000 2.635000 ;
      RECT  0.615000  0.805000  0.810000 0.970000 ;
      RECT  0.615000  0.970000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.245000 0.715000 ;
      RECT  1.020000  0.715000  1.245000 2.465000 ;
      RECT  1.435000  0.275000  1.805000 0.445000 ;
      RECT  1.435000  0.445000  1.605000 1.860000 ;
      RECT  1.435000  1.860000  3.250000 2.075000 ;
      RECT  1.435000  2.075000  1.710000 2.445000 ;
      RECT  1.880000  2.245000  2.210000 2.635000 ;
      RECT  1.975000  0.085000  2.305000 0.445000 ;
      RECT  2.120000  0.955000  2.465000 1.125000 ;
      RECT  2.120000  1.125000  2.290000 1.860000 ;
      RECT  2.695000  2.245000  3.590000 2.415000 ;
      RECT  2.820000  0.275000  3.595000 0.445000 ;
      RECT  3.080000  1.355000  3.275000 1.685000 ;
      RECT  3.080000  1.685000  3.250000 1.860000 ;
      RECT  3.420000  1.825000  4.385000 1.995000 ;
      RECT  3.420000  1.995000  3.590000 2.245000 ;
      RECT  3.425000  0.445000  3.595000 0.695000 ;
      RECT  3.425000  0.695000  4.385000 0.865000 ;
      RECT  3.760000  2.165000  3.930000 2.635000 ;
      RECT  3.765000  0.085000  3.965000 0.525000 ;
      RECT  4.215000  0.365000  4.565000 0.535000 ;
      RECT  4.215000  0.535000  4.385000 0.695000 ;
      RECT  4.215000  0.865000  4.385000 1.825000 ;
      RECT  4.215000  1.995000  4.385000 2.065000 ;
      RECT  4.215000  2.065000  4.450000 2.440000 ;
      RECT  4.555000  0.705000  5.135000 1.035000 ;
      RECT  4.555000  1.035000  4.795000 1.905000 ;
      RECT  4.695000  2.190000  5.765000 2.360000 ;
      RECT  4.735000  0.365000  5.475000 0.535000 ;
      RECT  4.985000  1.655000  5.425000 2.010000 ;
      RECT  5.305000  0.535000  5.475000 1.315000 ;
      RECT  5.305000  1.315000  6.105000 1.485000 ;
      RECT  5.595000  1.485000  6.105000 1.575000 ;
      RECT  5.595000  1.575000  5.765000 2.190000 ;
      RECT  5.645000  0.765000  6.445000 1.065000 ;
      RECT  5.645000  1.065000  5.815000 1.095000 ;
      RECT  5.725000  0.085000  6.095000 0.585000 ;
      RECT  5.935000  1.245000  6.105000 1.315000 ;
      RECT  5.935000  1.835000  6.105000 2.635000 ;
      RECT  6.275000  0.365000  6.735000 0.535000 ;
      RECT  6.275000  0.535000  6.445000 0.765000 ;
      RECT  6.275000  1.065000  6.445000 2.135000 ;
      RECT  6.275000  2.135000  6.525000 2.465000 ;
      RECT  6.615000  0.705000  7.165000 1.035000 ;
      RECT  6.615000  1.245000  6.805000 1.965000 ;
      RECT  6.750000  2.165000  7.635000 2.335000 ;
      RECT  6.965000  0.365000  7.505000 0.535000 ;
      RECT  6.975000  1.035000  7.165000 1.575000 ;
      RECT  6.975000  1.575000  7.295000 1.905000 ;
      RECT  7.335000  0.535000  7.505000 0.995000 ;
      RECT  7.335000  0.995000  8.400000 1.325000 ;
      RECT  7.335000  1.325000  7.635000 1.405000 ;
      RECT  7.465000  1.405000  7.635000 2.165000 ;
      RECT  7.750000  0.085000  8.120000 0.615000 ;
      RECT  7.805000  1.575000  8.755000 1.905000 ;
      RECT  7.815000  2.135000  8.120000 2.635000 ;
      RECT  8.390000  0.300000  8.750000 0.825000 ;
      RECT  8.470000  1.905000  8.755000 2.455000 ;
      RECT  8.570000  0.825000  8.750000 1.075000 ;
      RECT  8.570000  1.075000 10.485000 1.325000 ;
      RECT  8.570000  1.325000  8.755000 1.575000 ;
      RECT  8.925000  0.085000  9.095000 0.695000 ;
      RECT  8.925000  1.625000  9.105000 2.635000 ;
      RECT  9.795000  0.085000  9.965000 0.565000 ;
      RECT  9.795000  1.845000  9.965000 2.635000 ;
      RECT 10.635000  0.085000 10.805000 0.565000 ;
      RECT 10.635000  1.845000 10.805000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.615000  1.785000  0.785000 1.955000 ;
      RECT  1.055000  0.765000  1.225000 0.935000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.755000  0.765000  4.925000 0.935000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.215000  1.785000  5.385000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.625000  0.765000  6.795000 0.935000 ;
      RECT  6.625000  1.785000  6.795000 1.955000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.555000 1.755000 0.845000 1.800000 ;
      RECT 0.555000 1.800000 6.855000 1.940000 ;
      RECT 0.555000 1.940000 0.845000 1.985000 ;
      RECT 0.995000 0.735000 1.285000 0.780000 ;
      RECT 0.995000 0.780000 6.855000 0.920000 ;
      RECT 0.995000 0.920000 1.285000 0.965000 ;
      RECT 4.695000 0.735000 4.985000 0.780000 ;
      RECT 4.695000 0.920000 4.985000 0.965000 ;
      RECT 5.155000 1.755000 5.445000 1.800000 ;
      RECT 5.155000 1.940000 5.445000 1.985000 ;
      RECT 6.565000 0.735000 6.855000 0.780000 ;
      RECT 6.565000 0.920000 6.855000 0.965000 ;
      RECT 6.565000 1.755000 6.855000 1.800000 ;
      RECT 6.565000 1.940000 6.855000 1.985000 ;
  END
END sky130_fd_sc_hd__sdfxtp_4
MACRO sky130_fd_sc_hd__sdfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.460000 1.355000 2.790000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.260000 0.305000 9.605000 0.820000 ;
        RECT 9.260000 1.505000 9.605000 2.395000 ;
        RECT 9.435000 0.820000 9.605000 1.505000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.530000 1.035000 4.020000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.615000 3.250000 0.785000 ;
        RECT 1.780000 0.785000 1.950000 1.685000 ;
        RECT 2.475000 0.305000 2.650000 0.615000 ;
        RECT 3.080000 0.785000 3.250000 1.115000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.175000  0.345000  0.345000 0.635000 ;
      RECT 0.175000  0.635000  0.810000 0.805000 ;
      RECT 0.180000  1.795000  0.845000 1.965000 ;
      RECT 0.180000  1.965000  0.350000 2.465000 ;
      RECT 0.515000  0.085000  0.845000 0.465000 ;
      RECT 0.520000  2.135000  0.850000 2.635000 ;
      RECT 0.615000  0.805000  0.810000 0.970000 ;
      RECT 0.615000  0.970000  0.845000 1.795000 ;
      RECT 1.015000  0.345000  1.245000 0.715000 ;
      RECT 1.020000  0.715000  1.245000 2.465000 ;
      RECT 1.435000  0.275000  1.805000 0.445000 ;
      RECT 1.435000  0.445000  1.605000 1.860000 ;
      RECT 1.435000  1.860000  3.245000 2.075000 ;
      RECT 1.435000  2.075000  1.710000 2.445000 ;
      RECT 1.880000  2.245000  2.210000 2.635000 ;
      RECT 1.975000  0.085000  2.305000 0.445000 ;
      RECT 2.120000  0.955000  2.460000 1.125000 ;
      RECT 2.120000  1.125000  2.290000 1.860000 ;
      RECT 2.690000  2.245000  3.585000 2.415000 ;
      RECT 2.820000  0.275000  3.590000 0.445000 ;
      RECT 3.075000  1.355000  3.270000 1.685000 ;
      RECT 3.075000  1.685000  3.245000 1.860000 ;
      RECT 3.415000  1.825000  4.380000 1.995000 ;
      RECT 3.415000  1.995000  3.585000 2.245000 ;
      RECT 3.420000  0.445000  3.590000 0.695000 ;
      RECT 3.420000  0.695000  4.380000 0.865000 ;
      RECT 3.755000  2.165000  3.925000 2.635000 ;
      RECT 3.760000  0.085000  3.960000 0.525000 ;
      RECT 4.210000  0.365000  4.560000 0.535000 ;
      RECT 4.210000  0.535000  4.380000 0.695000 ;
      RECT 4.210000  0.865000  4.380000 1.825000 ;
      RECT 4.210000  1.995000  4.380000 2.065000 ;
      RECT 4.210000  2.065000  4.445000 2.440000 ;
      RECT 4.550000  0.705000  5.130000 1.035000 ;
      RECT 4.550000  1.035000  4.790000 1.905000 ;
      RECT 4.690000  2.190000  5.760000 2.360000 ;
      RECT 4.730000  0.365000  5.470000 0.535000 ;
      RECT 4.980000  1.655000  5.420000 2.010000 ;
      RECT 5.300000  0.535000  5.470000 1.315000 ;
      RECT 5.300000  1.315000  6.100000 1.485000 ;
      RECT 5.590000  1.485000  6.100000 1.575000 ;
      RECT 5.590000  1.575000  5.760000 2.190000 ;
      RECT 5.640000  0.765000  6.440000 1.065000 ;
      RECT 5.640000  1.065000  5.810000 1.095000 ;
      RECT 5.720000  0.085000  6.090000 0.585000 ;
      RECT 5.930000  1.245000  6.100000 1.315000 ;
      RECT 5.930000  1.835000  6.100000 2.635000 ;
      RECT 6.270000  0.365000  6.730000 0.535000 ;
      RECT 6.270000  0.535000  6.440000 0.765000 ;
      RECT 6.270000  1.065000  6.440000 2.135000 ;
      RECT 6.270000  2.135000  6.520000 2.465000 ;
      RECT 6.610000  0.705000  7.160000 1.035000 ;
      RECT 6.610000  1.245000  6.800000 1.965000 ;
      RECT 6.745000  2.165000  7.630000 2.335000 ;
      RECT 6.960000  0.365000  7.500000 0.535000 ;
      RECT 6.970000  1.035000  7.160000 1.575000 ;
      RECT 6.970000  1.575000  7.290000 1.905000 ;
      RECT 7.330000  0.535000  7.500000 0.995000 ;
      RECT 7.330000  0.995000  8.395000 1.325000 ;
      RECT 7.330000  1.325000  7.630000 1.405000 ;
      RECT 7.460000  1.405000  7.630000 2.165000 ;
      RECT 7.745000  0.085000  8.115000 0.615000 ;
      RECT 7.800000  1.575000  8.735000 1.905000 ;
      RECT 7.810000  2.135000  8.115000 2.635000 ;
      RECT 8.385000  0.300000  8.735000 0.825000 ;
      RECT 8.465000  1.905000  8.735000 2.455000 ;
      RECT 8.565000  0.825000  8.735000 0.995000 ;
      RECT 8.565000  0.995000  9.265000 1.325000 ;
      RECT 8.565000  1.325000  8.735000 1.575000 ;
      RECT 8.905000  0.085000  9.075000 0.695000 ;
      RECT 8.905000  1.625000  9.080000 2.635000 ;
      RECT 9.775000  0.085000  9.945000 0.930000 ;
      RECT 9.775000  1.405000  9.945000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.640000  1.785000 0.810000 1.955000 ;
      RECT 1.050000  0.765000 1.220000 0.935000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  0.765000 4.915000 0.935000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  1.785000 5.375000 1.955000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.620000  1.785000 6.790000 1.955000 ;
      RECT 6.630000  0.765000 6.800000 0.935000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 0.580000 1.755000 0.870000 1.800000 ;
      RECT 0.580000 1.800000 6.850000 1.940000 ;
      RECT 0.580000 1.940000 0.870000 1.985000 ;
      RECT 0.990000 0.735000 1.280000 0.780000 ;
      RECT 0.990000 0.780000 6.860000 0.920000 ;
      RECT 0.990000 0.920000 1.280000 0.965000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 6.560000 1.755000 6.850000 1.800000 ;
      RECT 6.560000 1.940000 6.850000 1.985000 ;
      RECT 6.570000 0.735000 6.860000 0.780000 ;
      RECT 6.570000 0.920000 6.860000 0.965000 ;
  END
END sky130_fd_sc_hd__sdfxtp_2
MACRO sky130_fd_sc_hd__sdfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.460000 1.355000 2.790000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.230000 0.305000 9.575000 0.820000 ;
        RECT 9.230000 1.505000 9.575000 2.395000 ;
        RECT 9.405000 0.820000 9.575000 1.505000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.530000 1.055000 3.990000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.760000 0.635000 3.250000 0.785000 ;
        RECT 1.760000 0.785000 1.990000 0.835000 ;
        RECT 1.760000 0.835000 1.930000 1.685000 ;
        RECT 1.870000 0.615000 3.250000 0.635000 ;
        RECT 2.475000 0.305000 2.650000 0.615000 ;
        RECT 3.065000 0.785000 3.250000 1.095000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.810000 0.805000 ;
      RECT 0.180000  1.795000 0.845000 1.965000 ;
      RECT 0.180000  1.965000 0.350000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.520000  2.135000 0.850000 2.635000 ;
      RECT 0.615000  0.805000 0.810000 0.970000 ;
      RECT 0.615000  0.970000 0.845000 1.795000 ;
      RECT 1.015000  0.345000 1.230000 0.715000 ;
      RECT 1.020000  0.715000 1.230000 2.465000 ;
      RECT 1.420000  0.260000 1.790000 0.465000 ;
      RECT 1.420000  0.465000 1.590000 1.860000 ;
      RECT 1.420000  1.860000 3.220000 2.075000 ;
      RECT 1.420000  2.075000 1.710000 2.445000 ;
      RECT 1.880000  2.245000 2.210000 2.635000 ;
      RECT 1.960000  0.085000 2.305000 0.445000 ;
      RECT 2.115000  0.960000 2.460000 1.130000 ;
      RECT 2.115000  1.130000 2.290000 1.860000 ;
      RECT 2.690000  2.245000 3.560000 2.415000 ;
      RECT 2.820000  0.275000 3.590000 0.445000 ;
      RECT 3.050000  1.305000 3.270000 1.635000 ;
      RECT 3.050000  1.635000 3.220000 1.860000 ;
      RECT 3.390000  1.825000 4.350000 1.995000 ;
      RECT 3.390000  1.995000 3.560000 2.245000 ;
      RECT 3.420000  0.445000 3.590000 0.715000 ;
      RECT 3.420000  0.715000 4.350000 0.885000 ;
      RECT 3.730000  2.165000 3.925000 2.635000 ;
      RECT 3.760000  0.085000 3.960000 0.545000 ;
      RECT 4.180000  0.285000 4.460000 0.615000 ;
      RECT 4.180000  0.615000 4.350000 0.715000 ;
      RECT 4.180000  0.885000 4.350000 1.825000 ;
      RECT 4.180000  1.995000 4.350000 2.065000 ;
      RECT 4.180000  2.065000 4.420000 2.440000 ;
      RECT 4.520000  0.780000 5.100000 1.035000 ;
      RECT 4.520000  1.035000 4.760000 1.905000 ;
      RECT 4.630000  0.705000 5.100000 0.780000 ;
      RECT 4.660000  2.190000 5.730000 2.360000 ;
      RECT 4.700000  0.365000 5.440000 0.535000 ;
      RECT 4.950000  1.655000 5.390000 2.010000 ;
      RECT 5.270000  0.535000 5.440000 1.315000 ;
      RECT 5.270000  1.315000 6.070000 1.485000 ;
      RECT 5.560000  1.485000 6.070000 1.575000 ;
      RECT 5.560000  1.575000 5.730000 2.190000 ;
      RECT 5.610000  0.765000 6.410000 1.065000 ;
      RECT 5.610000  1.065000 5.780000 1.095000 ;
      RECT 5.690000  0.085000 6.060000 0.585000 ;
      RECT 5.900000  1.245000 6.070000 1.315000 ;
      RECT 5.900000  1.835000 6.070000 2.635000 ;
      RECT 6.240000  0.365000 6.700000 0.535000 ;
      RECT 6.240000  0.535000 6.410000 0.765000 ;
      RECT 6.240000  1.065000 6.410000 2.135000 ;
      RECT 6.240000  2.135000 6.490000 2.465000 ;
      RECT 6.580000  0.705000 7.130000 1.035000 ;
      RECT 6.580000  1.245000 6.770000 1.965000 ;
      RECT 6.715000  2.165000 7.600000 2.335000 ;
      RECT 6.930000  0.365000 7.470000 0.535000 ;
      RECT 6.940000  1.035000 7.130000 1.575000 ;
      RECT 6.940000  1.575000 7.260000 1.905000 ;
      RECT 7.300000  0.535000 7.470000 0.995000 ;
      RECT 7.300000  0.995000 8.365000 1.325000 ;
      RECT 7.300000  1.325000 7.600000 1.405000 ;
      RECT 7.430000  1.405000 7.600000 2.165000 ;
      RECT 7.715000  0.085000 8.085000 0.615000 ;
      RECT 7.770000  1.575000 8.705000 1.905000 ;
      RECT 7.790000  2.135000 8.095000 2.635000 ;
      RECT 8.355000  0.300000 8.705000 0.825000 ;
      RECT 8.435000  1.905000 8.705000 2.455000 ;
      RECT 8.535000  0.825000 8.705000 0.995000 ;
      RECT 8.535000  0.995000 9.235000 1.325000 ;
      RECT 8.535000  1.325000 8.705000 1.575000 ;
      RECT 8.875000  0.085000 9.045000 0.695000 ;
      RECT 8.875000  1.625000 9.045000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.640000  1.785000 0.810000 1.955000 ;
      RECT 1.040000  0.765000 1.210000 0.935000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  0.765000 4.915000 0.935000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  1.785000 5.375000 1.955000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.590000  1.785000 6.760000 1.955000 ;
      RECT 6.630000  0.765000 6.800000 0.935000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
    LAYER met1 ;
      RECT 0.580000 1.755000 0.870000 1.800000 ;
      RECT 0.580000 1.800000 6.820000 1.940000 ;
      RECT 0.580000 1.940000 0.870000 1.985000 ;
      RECT 0.980000 0.735000 1.270000 0.780000 ;
      RECT 0.980000 0.780000 6.860000 0.920000 ;
      RECT 0.980000 0.920000 1.270000 0.965000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 6.530000 1.755000 6.820000 1.800000 ;
      RECT 6.530000 1.940000 6.820000 1.985000 ;
      RECT 6.570000 0.735000 6.860000 0.780000 ;
      RECT 6.570000 0.920000 6.860000 0.965000 ;
  END
END sky130_fd_sc_hd__sdfxtp_1
MACRO sky130_fd_sc_hd__bufbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufbuf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  5.235000 0.255000  5.485000 0.260000 ;
        RECT  5.235000 0.260000  5.565000 0.735000 ;
        RECT  5.235000 0.735000 11.875000 0.905000 ;
        RECT  5.235000 1.445000 11.875000 1.615000 ;
        RECT  5.235000 1.615000  5.565000 2.465000 ;
        RECT  6.075000 0.260000  6.405000 0.735000 ;
        RECT  6.075000 1.615000  6.405000 2.465000 ;
        RECT  6.155000 0.255000  6.325000 0.260000 ;
        RECT  6.915000 0.260000  7.245000 0.735000 ;
        RECT  6.915000 1.615000  7.245000 2.465000 ;
        RECT  6.995000 0.255000  7.165000 0.260000 ;
        RECT  7.755000 0.260000  8.085000 0.735000 ;
        RECT  7.755000 1.615000  8.085000 2.465000 ;
        RECT  8.595000 0.260000  8.925000 0.735000 ;
        RECT  8.595000 1.615000  8.925000 2.465000 ;
        RECT  9.435000 0.260000  9.765000 0.735000 ;
        RECT  9.435000 1.615000  9.765000 2.465000 ;
        RECT 10.275000 0.260000 10.605000 0.735000 ;
        RECT 10.275000 1.615000 10.605000 2.465000 ;
        RECT 11.115000 0.260000 11.445000 0.735000 ;
        RECT 11.115000 1.615000 11.445000 2.465000 ;
        RECT 11.620000 0.905000 11.875000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.175000  0.085000  0.345000 0.905000 ;
      RECT  0.175000  1.445000  0.345000 2.635000 ;
      RECT  0.515000  0.260000  0.845000 0.905000 ;
      RECT  0.515000  1.445000  0.845000 2.465000 ;
      RECT  0.610000  0.905000  0.845000 1.075000 ;
      RECT  0.610000  1.075000  2.205000 1.275000 ;
      RECT  0.610000  1.275000  0.845000 1.445000 ;
      RECT  1.035000  0.260000  1.365000 0.735000 ;
      RECT  1.035000  0.735000  2.545000 0.905000 ;
      RECT  1.035000  1.445000  2.545000 1.615000 ;
      RECT  1.035000  1.615000  1.365000 2.465000 ;
      RECT  1.535000  0.085000  1.705000 0.565000 ;
      RECT  1.535000  1.785000  1.705000 2.635000 ;
      RECT  1.875000  0.260000  2.205000 0.735000 ;
      RECT  1.875000  1.615000  2.205000 2.465000 ;
      RECT  2.375000  0.085000  2.545000 0.565000 ;
      RECT  2.375000  0.905000  2.545000 1.075000 ;
      RECT  2.375000  1.075000  4.685000 1.275000 ;
      RECT  2.375000  1.275000  2.545000 1.445000 ;
      RECT  2.375000  1.785000  2.545000 2.635000 ;
      RECT  2.715000  0.260000  3.045000 0.735000 ;
      RECT  2.715000  0.735000  5.065000 0.905000 ;
      RECT  2.715000  1.445000  5.065000 1.615000 ;
      RECT  2.715000  1.615000  3.045000 2.465000 ;
      RECT  3.215000  0.085000  3.385000 0.565000 ;
      RECT  3.215000  1.835000  3.385000 2.635000 ;
      RECT  3.555000  0.260000  3.885000 0.735000 ;
      RECT  3.555000  1.615000  3.885000 2.465000 ;
      RECT  4.055000  0.085000  4.225000 0.565000 ;
      RECT  4.055000  1.835000  4.225000 2.635000 ;
      RECT  4.395000  0.260000  4.725000 0.735000 ;
      RECT  4.395000  1.615000  4.725000 2.465000 ;
      RECT  4.890000  0.905000  5.065000 1.075000 ;
      RECT  4.890000  1.075000 11.450000 1.275000 ;
      RECT  4.890000  1.275000  5.065000 1.445000 ;
      RECT  4.895000  0.085000  5.065000 0.565000 ;
      RECT  4.895000  1.835000  5.065000 2.635000 ;
      RECT  5.735000  0.085000  5.905000 0.565000 ;
      RECT  5.735000  1.835000  5.905000 2.635000 ;
      RECT  6.575000  0.085000  6.745000 0.565000 ;
      RECT  6.575000  1.835000  6.745000 2.635000 ;
      RECT  7.415000  0.085000  7.585000 0.565000 ;
      RECT  7.415000  1.835000  7.585000 2.635000 ;
      RECT  8.255000  0.085000  8.425000 0.565000 ;
      RECT  8.255000  1.835000  8.425000 2.635000 ;
      RECT  9.095000  0.085000  9.265000 0.565000 ;
      RECT  9.095000  1.835000  9.265000 2.635000 ;
      RECT  9.935000  0.085000 10.105000 0.565000 ;
      RECT  9.935000  1.835000 10.105000 2.635000 ;
      RECT 10.775000  0.085000 10.945000 0.565000 ;
      RECT 10.775000  1.835000 10.945000 2.635000 ;
      RECT 11.615000  0.085000 11.785000 0.565000 ;
      RECT 11.615000  1.835000 11.785000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
  END
END sky130_fd_sc_hd__bufbuf_16
MACRO sky130_fd_sc_hd__bufbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufbuf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.230000 0.260000 3.560000 0.735000 ;
        RECT 3.230000 0.735000 6.815000 0.905000 ;
        RECT 3.230000 1.445000 6.815000 1.615000 ;
        RECT 3.230000 1.615000 3.560000 2.465000 ;
        RECT 4.070000 0.260000 4.400000 0.735000 ;
        RECT 4.070000 1.615000 4.400000 2.465000 ;
        RECT 4.910000 0.260000 5.240000 0.735000 ;
        RECT 4.910000 1.615000 5.240000 2.465000 ;
        RECT 5.750000 0.260000 6.080000 0.735000 ;
        RECT 5.750000 1.615000 6.080000 2.465000 ;
        RECT 6.435000 0.905000 6.815000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.095000  0.260000 0.425000 0.735000 ;
      RECT 0.095000  0.735000 0.780000 0.905000 ;
      RECT 0.095000  1.445000 0.780000 1.615000 ;
      RECT 0.095000  1.615000 0.425000 2.160000 ;
      RECT 0.595000  0.085000 0.765000 0.565000 ;
      RECT 0.595000  1.785000 0.765000 2.635000 ;
      RECT 0.610000  0.905000 0.780000 0.995000 ;
      RECT 0.610000  0.995000 1.040000 1.325000 ;
      RECT 0.610000  1.325000 0.780000 1.445000 ;
      RECT 1.000000  0.260000 1.380000 0.825000 ;
      RECT 1.000000  1.545000 1.380000 2.465000 ;
      RECT 1.210000  0.825000 1.380000 1.075000 ;
      RECT 1.210000  1.075000 2.720000 1.275000 ;
      RECT 1.210000  1.275000 1.380000 1.545000 ;
      RECT 1.550000  0.260000 1.880000 0.735000 ;
      RECT 1.550000  0.735000 3.060000 0.905000 ;
      RECT 1.550000  1.445000 3.060000 1.615000 ;
      RECT 1.550000  1.615000 1.880000 2.465000 ;
      RECT 2.050000  0.085000 2.220000 0.565000 ;
      RECT 2.050000  1.785000 2.220000 2.635000 ;
      RECT 2.390000  0.260000 2.720000 0.735000 ;
      RECT 2.390000  1.615000 2.720000 2.465000 ;
      RECT 2.890000  0.085000 3.060000 0.565000 ;
      RECT 2.890000  0.905000 3.060000 1.075000 ;
      RECT 2.890000  1.075000 5.360000 1.275000 ;
      RECT 2.890000  1.275000 3.060000 1.445000 ;
      RECT 2.890000  1.785000 3.060000 2.635000 ;
      RECT 3.730000  0.085000 3.900000 0.565000 ;
      RECT 3.730000  1.835000 3.900000 2.635000 ;
      RECT 4.570000  0.085000 4.740000 0.565000 ;
      RECT 4.570000  1.835000 4.740000 2.635000 ;
      RECT 5.410000  0.085000 5.580000 0.565000 ;
      RECT 5.410000  1.835000 5.580000 2.635000 ;
      RECT 6.250000  0.085000 6.420000 0.565000 ;
      RECT 6.250000  1.835000 6.420000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
END sky130_fd_sc_hd__bufbuf_8
MACRO sky130_fd_sc_hd__a2111oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.465000 0.985000 3.715000 1.445000 ;
        RECT 3.465000 1.445000 5.290000 1.675000 ;
        RECT 4.895000 0.995000 5.290000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.970000 1.015000 4.725000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.185000 1.030000 2.855000 1.275000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.045000 0.455000 1.445000 ;
        RECT 0.125000 1.445000 1.800000 1.680000 ;
        RECT 1.615000 1.030000 1.975000 1.275000 ;
        RECT 1.615000 1.275000 1.800000 1.445000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.755000 1.075000 1.425000 1.275000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.212750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.255000 0.380000 0.615000 ;
        RECT 0.120000 0.615000 5.355000 0.805000 ;
        RECT 0.120000 0.805000 3.255000 0.845000 ;
        RECT 0.900000 1.850000 2.140000 2.105000 ;
        RECT 1.050000 0.255000 1.295000 0.615000 ;
        RECT 1.965000 0.255000 2.295000 0.615000 ;
        RECT 1.970000 1.445000 3.255000 1.625000 ;
        RECT 1.970000 1.625000 2.140000 1.850000 ;
        RECT 2.965000 0.275000 3.295000 0.615000 ;
        RECT 3.025000 0.845000 3.255000 1.445000 ;
        RECT 5.020000 0.295000 5.355000 0.615000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.100000  1.870000 0.460000 2.275000 ;
      RECT 0.100000  2.275000 2.185000 2.295000 ;
      RECT 0.100000  2.295000 2.985000 2.465000 ;
      RECT 0.550000  0.085000 0.880000 0.445000 ;
      RECT 1.465000  0.085000 1.795000 0.445000 ;
      RECT 2.310000  1.795000 3.335000 1.845000 ;
      RECT 2.310000  1.845000 5.400000 1.965000 ;
      RECT 2.310000  1.965000 2.640000 2.060000 ;
      RECT 2.465000  0.085000 2.795000 0.445000 ;
      RECT 2.815000  2.135000 2.985000 2.295000 ;
      RECT 3.155000  1.965000 5.400000 2.095000 ;
      RECT 3.155000  2.095000 3.520000 2.465000 ;
      RECT 3.690000  2.275000 4.020000 2.635000 ;
      RECT 4.125000  0.085000 4.455000 0.445000 ;
      RECT 4.190000  2.095000 5.400000 2.105000 ;
      RECT 4.190000  2.105000 4.400000 2.465000 ;
      RECT 4.570000  2.275000 4.900000 2.635000 ;
      RECT 5.070000  2.105000 5.400000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111oi_2
MACRO sky130_fd_sc_hd__a2111oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095000 1.020000 7.745000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.960000 1.020000 9.990000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.955000 1.020000 5.650000 1.275000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055000 1.020000 3.745000 1.275000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495000 1.020000 1.845000 1.275000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  2.009500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.615000 7.620000 0.785000 ;
        RECT 0.145000 0.785000 0.320000 1.475000 ;
        RECT 0.145000 1.475000 1.720000 1.655000 ;
        RECT 0.530000 1.655000 1.720000 1.685000 ;
        RECT 0.530000 1.685000 0.860000 2.085000 ;
        RECT 0.615000 0.455000 0.790000 0.615000 ;
        RECT 1.390000 1.685000 1.720000 2.085000 ;
        RECT 1.460000 0.455000 1.650000 0.615000 ;
        RECT 2.400000 0.455000 2.590000 0.615000 ;
        RECT 3.260000 0.455000 3.510000 0.615000 ;
        RECT 4.180000 0.455000 4.420000 0.615000 ;
        RECT 5.090000 0.455000 5.275000 0.615000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.100000  1.835000  0.360000 2.255000 ;
      RECT 0.100000  2.255000  3.870000 2.445000 ;
      RECT 0.115000  0.085000  0.445000 0.445000 ;
      RECT 0.960000  0.085000  1.290000 0.445000 ;
      RECT 1.030000  1.855000  1.220000 2.255000 ;
      RECT 1.820000  0.085000  2.230000 0.445000 ;
      RECT 1.890000  1.855000  2.080000 2.255000 ;
      RECT 2.250000  1.475000  5.680000 1.655000 ;
      RECT 2.250000  1.655000  3.440000 1.685000 ;
      RECT 2.250000  1.685000  2.580000 2.085000 ;
      RECT 2.750000  1.855000  2.940000 2.255000 ;
      RECT 2.760000  0.085000  3.090000 0.445000 ;
      RECT 3.110000  1.685000  3.440000 2.085000 ;
      RECT 3.610000  1.835000  3.870000 2.255000 ;
      RECT 3.680000  0.085000  4.010000 0.445000 ;
      RECT 4.060000  1.835000  4.320000 2.255000 ;
      RECT 4.060000  2.255000  5.180000 2.275000 ;
      RECT 4.060000  2.275000  6.050000 2.445000 ;
      RECT 4.490000  1.655000  5.680000 1.685000 ;
      RECT 4.490000  1.685000  4.820000 2.085000 ;
      RECT 4.590000  0.085000  4.920000 0.445000 ;
      RECT 4.990000  1.855000  5.180000 2.255000 ;
      RECT 5.350000  1.685000  5.680000 2.085000 ;
      RECT 5.445000  0.085000  5.780000 0.445000 ;
      RECT 5.860000  1.445000  9.770000 1.615000 ;
      RECT 5.860000  1.615000  6.050000 2.275000 ;
      RECT 5.980000  0.275000  8.075000 0.445000 ;
      RECT 6.220000  1.785000  6.550000 2.635000 ;
      RECT 6.720000  1.615000  6.910000 2.315000 ;
      RECT 7.080000  1.805000  7.410000 2.635000 ;
      RECT 7.580000  1.615000  9.770000 1.665000 ;
      RECT 7.580000  1.665000  7.910000 2.315000 ;
      RECT 7.885000  0.445000  8.075000 0.615000 ;
      RECT 7.885000  0.615000  9.865000 0.785000 ;
      RECT 8.080000  1.895000  8.410000 2.635000 ;
      RECT 8.245000  0.085000  8.575000 0.445000 ;
      RECT 8.580000  1.665000  9.770000 1.670000 ;
      RECT 8.580000  1.670000  8.840000 2.290000 ;
      RECT 8.745000  0.300000  8.935000 0.615000 ;
      RECT 9.030000  1.915000  9.360000 2.635000 ;
      RECT 9.105000  0.085000  9.435000 0.445000 ;
      RECT 9.530000  1.670000  9.770000 2.260000 ;
      RECT 9.605000  0.290000  9.865000 0.615000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111oi_4
MACRO sky130_fd_sc_hd__a2111oi_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035000 1.070000 2.625000 1.400000 ;
        RECT 2.355000 0.660000 2.625000 1.070000 ;
        RECT 2.355000 1.400000 2.625000 1.735000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.795000 0.650000 3.135000 1.735000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 1.055000 1.845000 1.735000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.055000 1.325000 2.360000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.730000 0.435000 1.655000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  0.424000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.825000 0.785000 2.465000 ;
        RECT 0.605000 0.635000 2.040000 0.885000 ;
        RECT 0.605000 0.885000 0.785000 1.825000 ;
        RECT 0.785000 0.255000 1.040000 0.615000 ;
        RECT 0.785000 0.615000 2.040000 0.635000 ;
        RECT 1.710000 0.280000 2.040000 0.615000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.285000  0.085000 0.615000 0.465000 ;
      RECT 1.210000  0.085000 1.540000 0.445000 ;
      RECT 1.540000  1.905000 2.870000 2.085000 ;
      RECT 1.540000  2.085000 1.870000 2.465000 ;
      RECT 2.040000  2.255000 2.370000 2.635000 ;
      RECT 2.470000  0.085000 2.800000 0.480000 ;
      RECT 2.540000  2.085000 2.870000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111oi_0
MACRO sky130_fd_sc_hd__a2111oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 0.995000 2.725000 1.400000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.350000 3.090000 1.020000 ;
        RECT 2.905000 1.020000 3.540000 1.290000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 1.050000 2.270000 1.400000 ;
        RECT 1.940000 1.400000 2.215000 2.455000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 1.050000 1.770000 2.455000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.785000 1.050000 1.235000 2.455000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.388750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.700000 1.375000 0.705000 ;
        RECT 0.145000 0.705000 2.420000 0.815000 ;
        RECT 0.145000 0.815000 2.300000 0.880000 ;
        RECT 0.145000 0.880000 0.530000 2.460000 ;
        RECT 1.045000 0.260000 1.375000 0.700000 ;
        RECT 2.090000 0.305000 2.420000 0.705000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
    PORT
      LAYER pwell ;
        RECT 1.975000 -0.065000 2.145000 0.105000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.315000  0.085000 0.630000 0.525000 ;
      RECT 1.550000  0.085000 1.880000 0.535000 ;
      RECT 2.395000  1.580000 3.505000 1.750000 ;
      RECT 2.395000  1.750000 2.625000 2.460000 ;
      RECT 2.800000  1.920000 3.130000 2.635000 ;
      RECT 3.270000  0.085000 3.510000 0.760000 ;
      RECT 3.310000  1.750000 3.505000 2.460000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111oi_1
MACRO sky130_fd_sc_hd__a211oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655000 1.075000 3.005000 1.245000 ;
        RECT 1.660000 1.035000 3.005000 1.075000 ;
        RECT 1.660000 1.245000 3.005000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.035000 1.385000 1.445000 ;
        RECT 0.100000 1.445000 3.575000 1.625000 ;
        RECT 3.245000 1.035000 3.575000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.745000 1.035000 4.755000 1.275000 ;
        RECT 3.745000 1.275000 4.460000 1.615000 ;
      LAYER mcon ;
        RECT 3.830000 1.445000 4.000000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.590000 0.995000 6.935000 1.325000 ;
        RECT 6.590000 1.325000 6.760000 1.615000 ;
      LAYER mcon ;
        RECT 6.590000 1.445000 6.760000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.770000 1.415000 4.060000 1.460000 ;
        RECT 3.770000 1.460000 6.820000 1.600000 ;
        RECT 3.770000 1.600000 4.060000 1.645000 ;
        RECT 6.530000 1.415000 6.820000 1.460000 ;
        RECT 6.530000 1.600000 6.820000 1.645000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.000000 1.035000 6.350000 1.275000 ;
        RECT 6.130000 1.275000 6.350000 1.695000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.685000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775000 0.675000 3.330000 0.695000 ;
        RECT 1.775000 0.695000 7.275000 0.825000 ;
        RECT 1.775000 0.825000 6.355000 0.865000 ;
        RECT 3.875000 0.255000 4.195000 0.615000 ;
        RECT 3.875000 0.615000 5.045000 0.625000 ;
        RECT 3.875000 0.625000 7.275000 0.695000 ;
        RECT 4.875000 0.255000 5.045000 0.615000 ;
        RECT 5.170000 1.865000 7.275000 2.085000 ;
        RECT 5.715000 0.255000 5.885000 0.615000 ;
        RECT 5.715000 0.615000 7.275000 0.625000 ;
        RECT 6.930000 1.495000 7.275000 1.865000 ;
        RECT 7.105000 0.825000 7.275000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.095000  0.085000 0.395000 0.585000 ;
      RECT 0.095000  1.795000 3.705000 2.085000 ;
      RECT 0.095000  2.085000 0.345000 2.465000 ;
      RECT 0.515000  2.255000 0.845000 2.635000 ;
      RECT 0.565000  0.530000 0.775000 0.695000 ;
      RECT 0.565000  0.695000 1.605000 0.865000 ;
      RECT 0.950000  0.085000 1.185000 0.525000 ;
      RECT 1.015000  2.085000 3.705000 2.105000 ;
      RECT 1.015000  2.105000 1.185000 2.465000 ;
      RECT 1.355000  0.255000 3.365000 0.505000 ;
      RECT 1.355000  0.505000 1.605000 0.695000 ;
      RECT 1.355000  2.275000 1.685000 2.635000 ;
      RECT 1.855000  2.105000 2.025000 2.465000 ;
      RECT 2.195000  2.275000 2.525000 2.635000 ;
      RECT 2.695000  2.105000 2.865000 2.465000 ;
      RECT 3.035000  2.275000 3.365000 2.635000 ;
      RECT 3.535000  0.085000 3.705000 0.525000 ;
      RECT 3.535000  2.105000 3.705000 2.255000 ;
      RECT 3.535000  2.255000 7.270000 2.465000 ;
      RECT 3.875000  1.785000 4.910000 2.085000 ;
      RECT 4.365000  0.085000 4.695000 0.445000 ;
      RECT 4.630000  1.445000 5.960000 1.695000 ;
      RECT 4.630000  1.695000 4.910000 1.785000 ;
      RECT 5.215000  0.085000 5.545000 0.445000 ;
      RECT 6.055000  0.085000 6.385000 0.445000 ;
      RECT 6.915000  0.085000 7.270000 0.445000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__a211oi_4
MACRO sky130_fd_sc_hd__a211oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.265000 0.855000 0.995000 ;
        RECT 0.605000 0.995000 1.245000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.765000 0.435000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.425000 0.995000 1.755000 1.325000 ;
        RECT 1.525000 1.325000 1.755000 2.455000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.995000 2.235000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.619250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.180000 0.265000 1.365000 0.625000 ;
        RECT 1.180000 0.625000 2.660000 0.815000 ;
        RECT 1.935000 1.785000 2.660000 2.455000 ;
        RECT 2.055000 0.265000 2.280000 0.625000 ;
        RECT 2.445000 0.815000 2.660000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  0.085000 0.425000 0.595000 ;
      RECT 0.250000  1.525000 1.355000 1.725000 ;
      RECT 0.250000  1.725000 0.500000 2.455000 ;
      RECT 0.670000  1.905000 1.000000 2.635000 ;
      RECT 1.170000  1.725000 1.355000 2.455000 ;
      RECT 1.545000  0.085000 1.875000 0.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__a211oi_1
MACRO sky130_fd_sc_hd__a211oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.370000 1.035000 3.080000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.740000 1.035000 4.500000 1.285000 ;
        RECT 4.175000 1.285000 4.500000 1.655000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.035000 1.785000 1.285000 ;
        RECT 1.035000 1.285000 1.255000 1.615000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.995000 0.405000 1.615000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.826000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 0.255000 0.835000 0.655000 ;
        RECT 0.575000 0.655000 3.145000 0.855000 ;
        RECT 0.575000 0.855000 0.855000 1.785000 ;
        RECT 0.575000 1.785000 0.905000 2.105000 ;
        RECT 1.505000 0.285000 1.695000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.125000 -0.085000 0.295000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.145000  0.085000 0.395000 0.815000 ;
      RECT 0.145000  1.785000 0.405000 2.285000 ;
      RECT 0.145000  2.285000 2.215000 2.455000 ;
      RECT 1.005000  0.085000 1.335000 0.475000 ;
      RECT 1.075000  1.785000 1.265000 2.255000 ;
      RECT 1.075000  2.255000 2.215000 2.285000 ;
      RECT 1.435000  1.455000 3.975000 1.655000 ;
      RECT 1.435000  1.655000 1.765000 2.075000 ;
      RECT 1.865000  0.085000 2.195000 0.475000 ;
      RECT 1.935000  1.835000 2.215000 2.255000 ;
      RECT 2.385000  0.265000 3.495000 0.475000 ;
      RECT 2.435000  1.835000 2.665000 2.635000 ;
      RECT 2.845000  1.655000 3.115000 2.465000 ;
      RECT 3.295000  1.835000 3.525000 2.635000 ;
      RECT 3.325000  0.475000 3.495000 0.635000 ;
      RECT 3.325000  0.635000 4.435000 0.855000 ;
      RECT 3.675000  0.085000 4.005000 0.455000 ;
      RECT 3.705000  1.655000 3.975000 2.465000 ;
      RECT 4.155000  1.835000 4.385000 2.635000 ;
      RECT 4.185000  0.265000 4.435000 0.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__a211oi_2
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.402500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.290000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 2.370000 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 6.170000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 6.440000 5.680000 ;
      LAYER pwell ;
        RECT 0.145000 4.595000 0.315000 5.120000 ;
        RECT 5.925000 4.595000 6.095000 5.120000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.500000 6.170000 3.640000 ;
        RECT 0.080000 3.455000 0.370000 3.500000 ;
        RECT 0.080000 3.640000 0.370000 3.685000 ;
        RECT 5.870000 3.455000 6.160000 3.500000 ;
        RECT 5.870000 3.640000 6.160000 3.685000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 4.135000 ;
        RECT  4.250000 1.305000 6.630000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 6.440000 5.525000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  2.985000 0.375000 3.970000 ;
      RECT 0.085000  4.630000 0.375000 5.355000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.290000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.290000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 6.440000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.865000  0.085000 6.155000 0.810000 ;
      RECT 5.865000  2.985000 6.155000 3.955000 ;
      RECT 5.865000  4.630000 6.155000 5.355000 ;
    LAYER mcon ;
      RECT 0.140000  3.485000 0.310000 3.655000 ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 5.930000  3.485000 6.100000 3.655000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 6.440000 0.240000 ;
    LAYER pwell ;
      RECT 0.145000 0.320000 0.315000 0.845000 ;
      RECT 5.925000 0.320000 6.095000 0.845000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.072500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.255000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 1.085000 ;
        RECT 5.360000 1.085000 6.555000 1.410000 ;
        RECT 5.360000 1.410000 5.635000 2.370000 ;
        RECT 6.280000 1.410000 6.555000 2.370000 ;
        RECT 6.335000 0.255000 6.555000 1.085000 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 7.290000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 7.360000 5.680000 ;
      LAYER pwell ;
        RECT 0.145000 4.595000 0.315000 5.120000 ;
        RECT 7.045000 4.595000 7.215000 5.120000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.500000 7.290000 3.640000 ;
        RECT 0.080000 3.455000 0.370000 3.500000 ;
        RECT 0.080000 3.640000 0.370000 3.685000 ;
        RECT 6.930000 3.455000 7.220000 3.500000 ;
        RECT 6.930000 3.640000 7.220000 3.685000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 4.135000 ;
        RECT  4.250000 1.305000 7.405000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 7.360000 5.525000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  2.985000 0.375000 3.970000 ;
      RECT 0.085000  4.630000 0.375000 5.355000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.255000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.255000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 7.360000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.825000  0.085000 6.155000 0.845000 ;
      RECT 5.905000  1.610000 6.075000 2.635000 ;
      RECT 6.755000  0.085000 7.005000 0.925000 ;
      RECT 6.755000  1.610000 6.935000 2.635000 ;
      RECT 6.985000  2.985000 7.275000 3.955000 ;
      RECT 6.985000  4.630000 7.275000 5.355000 ;
    LAYER mcon ;
      RECT 0.140000  3.485000 0.310000 3.655000 ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.585000  5.355000 6.755000 5.525000 ;
      RECT 6.990000  3.485000 7.160000 3.655000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.045000  5.355000 7.215000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 7.360000 0.240000 ;
    LAYER pwell ;
      RECT 0.145000 0.320000 0.315000 0.845000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.070000 3.290000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.610500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335000 0.255000 5.635000 0.980000 ;
        RECT 5.360000 0.980000 5.635000 2.370000 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.380000 2.065000 2.390000 2.335000 ;
        RECT 2.060000 1.635000 2.390000 2.065000 ;
        RECT 2.060000 2.335000 2.390000 2.660000 ;
        RECT 2.060000 2.660000 2.810000 3.750000 ;
      LAYER mcon ;
        RECT 1.420000 2.115000 1.590000 2.285000 ;
        RECT 1.780000 2.115000 1.950000 2.285000 ;
        RECT 2.140000 2.115000 2.310000 2.285000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 2.140000 6.370000 2.280000 ;
        RECT 1.360000 2.085000 2.370000 2.140000 ;
        RECT 1.360000 2.280000 2.370000 2.315000 ;
      LAYER nwell ;
        RECT 1.920000 1.305000 2.980000 4.135000 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 6.440000 5.680000 ;
      LAYER pwell ;
        RECT 0.145000 4.595000 0.315000 5.120000 ;
        RECT 6.125000 4.595000 6.295000 5.120000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.500000 6.300000 3.640000 ;
        RECT 0.080000 3.455000 0.370000 3.500000 ;
        RECT 0.080000 3.640000 0.370000 3.685000 ;
        RECT 6.010000 3.455000 6.300000 3.500000 ;
        RECT 6.010000 3.640000 6.300000 3.685000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 4.135000 ;
        RECT  4.250000 1.305000 6.630000 4.135000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 1.890000 2.805000 ;
      RECT 0.000000  5.355000 6.440000 5.525000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  2.985000 0.375000 3.970000 ;
      RECT 0.085000  4.630000 0.375000 5.355000 ;
      RECT 2.020000  0.085000 2.350000 0.895000 ;
      RECT 2.560000  0.375000 2.800000 2.130000 ;
      RECT 2.560000  2.130000 3.390000 2.370000 ;
      RECT 2.645000  4.515000 2.905000 5.355000 ;
      RECT 3.060000  2.370000 3.390000 3.965000 ;
      RECT 3.075000  4.265000 4.265000 4.325000 ;
      RECT 3.075000  4.325000 3.405000 5.185000 ;
      RECT 3.115000  0.085000 3.445000 0.900000 ;
      RECT 3.145000  4.155000 4.195000 4.265000 ;
      RECT 3.575000  4.515000 3.765000 5.355000 ;
      RECT 3.615000  0.255000 3.805000 0.730000 ;
      RECT 3.615000  0.730000 4.665000 0.980000 ;
      RECT 3.680000  2.405000 4.190000 2.575000 ;
      RECT 3.680000  2.575000 3.850000 3.470000 ;
      RECT 3.680000  3.470000 4.720000 3.640000 ;
      RECT 3.935000  4.325000 4.265000 5.185000 ;
      RECT 3.975000  0.085000 4.305000 0.560000 ;
      RECT 4.020000  0.980000 4.190000 2.405000 ;
      RECT 4.020000  2.745000 4.640000 2.915000 ;
      RECT 4.020000  2.915000 4.190000 3.300000 ;
      RECT 4.020000  3.810000 4.190000 4.155000 ;
      RECT 4.390000  3.085000 4.720000 3.470000 ;
      RECT 4.410000  3.640000 4.720000 3.740000 ;
      RECT 4.445000  4.515000 4.955000 5.355000 ;
      RECT 4.470000  1.625000 4.640000 2.745000 ;
      RECT 4.475000  0.255000 4.665000 0.730000 ;
      RECT 4.835000  0.085000 5.165000 0.900000 ;
      RECT 4.890000  1.625000 5.120000 2.635000 ;
      RECT 4.890000  2.635000 6.440000 2.805000 ;
      RECT 4.890000  2.805000 5.120000 3.740000 ;
      RECT 5.135000  4.405000 5.765000 4.460000 ;
      RECT 5.135000  4.460000 5.695000 4.820000 ;
      RECT 5.135000  4.820000 5.485000 5.160000 ;
      RECT 5.360000  3.070000 5.550000 4.125000 ;
      RECT 5.360000  4.125000 6.085000 4.355000 ;
      RECT 5.360000  4.355000 5.765000 4.405000 ;
      RECT 5.825000  0.085000 6.155000 0.900000 ;
      RECT 5.905000  1.610000 6.075000 2.635000 ;
      RECT 6.065000  2.985000 6.355000 3.955000 ;
      RECT 6.065000  4.630000 6.355000 5.355000 ;
    LAYER mcon ;
      RECT 0.140000  3.485000 0.310000 3.655000 ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.145000  5.355000 0.315000 5.525000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.605000  5.355000 0.775000 5.525000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.065000  5.355000 1.235000 5.525000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.525000  5.355000 1.695000 5.525000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  5.355000 2.155000 5.525000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  5.355000 2.615000 5.525000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  5.355000 3.075000 5.525000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  5.355000 3.535000 5.525000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  5.355000 3.995000 5.525000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  5.355000 4.455000 5.525000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  5.355000 4.915000 5.525000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.205000  5.355000 5.375000 5.525000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.665000  5.355000 5.835000 5.525000 ;
      RECT 6.070000  3.485000 6.240000 3.655000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.125000  5.355000 6.295000 5.525000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 6.440000 0.240000 ;
    LAYER pwell ;
      RECT 0.145000 0.320000 0.315000 0.845000 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2
MACRO sky130_fd_sc_hd__edfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__edfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.465000 0.305000 10.795000 2.420000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.795000  1.125000  4.980000 1.720000 ;
      RECT  4.815000  0.735000  5.320000 0.955000 ;
      RECT  4.915000  2.175000  5.955000 2.375000 ;
      RECT  5.005000  0.255000  5.680000 0.565000 ;
      RECT  5.150000  0.955000  5.320000 1.655000 ;
      RECT  5.150000  1.655000  5.615000 2.005000 ;
      RECT  5.510000  0.565000  5.680000 1.315000 ;
      RECT  5.510000  1.315000  6.360000 1.485000 ;
      RECT  5.785000  1.485000  6.360000 1.575000 ;
      RECT  5.785000  1.575000  5.955000 2.175000 ;
      RECT  5.870000  0.765000  6.935000 1.045000 ;
      RECT  5.870000  1.045000  7.445000 1.065000 ;
      RECT  5.870000  1.065000  6.070000 1.095000 ;
      RECT  5.945000  0.085000  6.340000 0.560000 ;
      RECT  6.125000  1.835000  6.360000 2.635000 ;
      RECT  6.190000  1.245000  6.360000 1.315000 ;
      RECT  6.530000  0.255000  6.935000 0.765000 ;
      RECT  6.530000  1.065000  7.445000 1.375000 ;
      RECT  6.530000  1.375000  6.860000 2.465000 ;
      RECT  7.070000  2.105000  7.360000 2.635000 ;
      RECT  7.165000  0.085000  7.440000 0.615000 ;
      RECT  7.790000  1.245000  7.980000 1.965000 ;
      RECT  7.925000  2.165000  8.810000 2.355000 ;
      RECT  8.005000  0.705000  8.470000 1.035000 ;
      RECT  8.025000  0.330000  8.810000 0.535000 ;
      RECT  8.150000  1.035000  8.470000 1.995000 ;
      RECT  8.640000  0.535000  8.810000 0.995000 ;
      RECT  8.640000  0.995000  9.510000 1.325000 ;
      RECT  8.640000  1.325000  8.810000 2.165000 ;
      RECT  8.980000  1.530000  9.880000 1.905000 ;
      RECT  8.980000  2.135000  9.240000 2.635000 ;
      RECT  9.050000  0.085000  9.365000 0.615000 ;
      RECT  9.540000  1.905000  9.880000 2.465000 ;
      RECT  9.550000  0.300000  9.880000 0.825000 ;
      RECT  9.690000  0.825000  9.880000 1.530000 ;
      RECT 10.050000  0.085000 10.295000 0.900000 ;
      RECT 10.050000  1.465000 10.295000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.800000  1.445000  4.970000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.210000  1.785000  5.380000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.800000  1.785000  7.970000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.220000  1.445000  8.390000 1.615000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.700000  0.765000  9.870000 0.935000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.575000 1.755000 0.865000 1.800000 ;
      RECT 0.575000 1.800000 8.030000 1.940000 ;
      RECT 0.575000 1.940000 0.865000 1.985000 ;
      RECT 0.955000 1.415000 1.245000 1.460000 ;
      RECT 0.955000 1.460000 8.450000 1.600000 ;
      RECT 0.955000 1.600000 1.245000 1.645000 ;
      RECT 1.295000 0.395000 4.415000 0.580000 ;
      RECT 1.295000 0.580000 1.585000 0.625000 ;
      RECT 3.745000 0.735000 4.035000 0.780000 ;
      RECT 3.745000 0.780000 9.930000 0.920000 ;
      RECT 3.745000 0.920000 4.035000 0.965000 ;
      RECT 4.125000 0.580000 4.415000 0.625000 ;
      RECT 4.740000 1.415000 5.030000 1.460000 ;
      RECT 4.740000 1.600000 5.030000 1.645000 ;
      RECT 5.150000 1.755000 5.440000 1.800000 ;
      RECT 5.150000 1.940000 5.440000 1.985000 ;
      RECT 7.740000 1.755000 8.030000 1.800000 ;
      RECT 7.740000 1.940000 8.030000 1.985000 ;
      RECT 8.160000 1.415000 8.450000 1.460000 ;
      RECT 8.160000 1.600000 8.450000 1.645000 ;
      RECT 9.640000 0.735000 9.930000 0.780000 ;
      RECT 9.640000 0.920000 9.930000 0.965000 ;
  END
END sky130_fd_sc_hd__edfxtp_1
MACRO sky130_fd_sc_hd__fa_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fa_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.631500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245000 0.995000 1.755000 1.275000 ;
        RECT 1.245000 1.275000 1.505000 1.325000 ;
      LAYER mcon ;
        RECT 1.525000 1.105000 1.695000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.685000 1.030000 3.075000 1.360000 ;
      LAYER mcon ;
        RECT 2.905000 1.105000 3.075000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.720000 0.955000 5.080000 1.275000 ;
      LAYER mcon ;
        RECT 4.765000 1.105000 4.935000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.105000 0.995000 6.960000 1.275000 ;
      LAYER mcon ;
        RECT 6.145000 1.105000 6.315000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465000 1.075000 1.755000 1.120000 ;
        RECT 1.465000 1.120000 6.375000 1.260000 ;
        RECT 1.465000 1.260000 1.755000 1.305000 ;
        RECT 2.845000 1.075000 3.135000 1.120000 ;
        RECT 2.845000 1.260000 3.135000 1.305000 ;
        RECT 4.705000 1.075000 4.995000 1.120000 ;
        RECT 4.705000 1.260000 4.995000 1.305000 ;
        RECT 6.085000 1.075000 6.375000 1.120000 ;
        RECT 6.085000 1.260000 6.375000 1.305000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.631500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.645000 1.445000 2.155000 1.690000 ;
      LAYER mcon ;
        RECT 1.985000 1.445000 2.155000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.655000 1.435000 4.070000 1.745000 ;
      LAYER mcon ;
        RECT 3.845000 1.445000 4.015000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.150000 1.445000 6.835000 1.735000 ;
      LAYER mcon ;
        RECT 6.605000 1.445000 6.775000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.925000 1.415000 2.215000 1.460000 ;
        RECT 1.925000 1.460000 6.835000 1.600000 ;
        RECT 1.925000 1.600000 2.215000 1.645000 ;
        RECT 3.785000 1.415000 4.075000 1.460000 ;
        RECT 3.785000 1.600000 4.075000 1.645000 ;
        RECT 6.545000 1.415000 6.835000 1.460000 ;
        RECT 6.545000 1.600000 6.835000 1.645000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.475500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.125000 1.105000 2.495000 1.275000 ;
        RECT 2.325000 1.275000 2.495000 1.570000 ;
        RECT 2.325000 1.570000 3.415000 1.740000 ;
        RECT 3.245000 0.965000 4.465000 1.250000 ;
        RECT 3.245000 1.250000 3.415000 1.570000 ;
        RECT 4.295000 1.250000 4.465000 1.435000 ;
        RECT 4.295000 1.435000 4.655000 1.515000 ;
        RECT 4.295000 1.515000 5.920000 1.685000 ;
        RECT 5.670000 1.355000 5.920000 1.515000 ;
        RECT 5.670000 1.685000 5.920000 1.955000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.735000 0.690000 0.905000 ;
        RECT 0.085000 0.905000 0.370000 1.415000 ;
        RECT 0.085000 1.415000 0.735000 1.585000 ;
        RECT 0.520000 0.315000 0.850000 0.485000 ;
        RECT 0.520000 0.485000 0.690000 0.735000 ;
        RECT 0.565000 1.585000 0.735000 1.780000 ;
        RECT 0.565000 1.780000 0.810000 1.950000 ;
        RECT 0.600000 1.950000 0.810000 2.465000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.523500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.395000 0.255000 7.725000 0.485000 ;
        RECT 7.395000 1.795000 7.645000 1.965000 ;
        RECT 7.395000 1.965000 7.565000 2.465000 ;
        RECT 7.475000 0.485000 7.725000 0.735000 ;
        RECT 7.475000 0.735000 8.195000 0.905000 ;
        RECT 7.475000 1.415000 8.195000 1.585000 ;
        RECT 7.475000 1.585000 7.645000 1.795000 ;
        RECT 7.970000 0.905000 8.195000 1.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.180000  0.085000 0.350000 0.565000 ;
      RECT 0.180000  1.795000 0.350000 2.635000 ;
      RECT 0.540000  1.075000 1.075000 1.245000 ;
      RECT 0.905000  0.655000 2.165000 0.825000 ;
      RECT 0.905000  0.825000 1.075000 1.075000 ;
      RECT 0.905000  1.245000 1.075000 1.430000 ;
      RECT 0.905000  1.430000 1.110000 1.495000 ;
      RECT 0.905000  1.495000 1.475000 1.600000 ;
      RECT 0.940000  1.600000 1.475000 1.665000 ;
      RECT 0.980000  2.275000 1.310000 2.635000 ;
      RECT 1.020000  0.085000 1.350000 0.465000 ;
      RECT 1.305000  1.665000 1.475000 1.910000 ;
      RECT 1.305000  1.910000 2.245000 2.080000 ;
      RECT 1.535000  0.255000 2.165000 0.655000 ;
      RECT 1.900000  2.080000 2.245000 2.465000 ;
      RECT 1.925000  0.825000 2.165000 0.935000 ;
      RECT 2.415000  0.255000 2.585000 0.615000 ;
      RECT 2.415000  0.615000 3.425000 0.785000 ;
      RECT 2.415000  1.935000 3.490000 2.105000 ;
      RECT 2.415000  2.105000 2.585000 2.465000 ;
      RECT 2.755000  0.085000 3.085000 0.445000 ;
      RECT 2.755000  2.275000 3.085000 2.635000 ;
      RECT 3.255000  0.255000 3.425000 0.615000 ;
      RECT 3.255000  2.105000 3.490000 2.465000 ;
      RECT 3.695000  0.085000 4.025000 0.490000 ;
      RECT 3.695000  1.915000 4.025000 2.635000 ;
      RECT 4.195000  0.255000 4.365000 0.615000 ;
      RECT 4.195000  0.615000 5.205000 0.785000 ;
      RECT 4.195000  1.935000 5.205000 2.105000 ;
      RECT 4.195000  2.105000 4.365000 2.465000 ;
      RECT 4.535000  0.085000 4.865000 0.445000 ;
      RECT 4.535000  2.275000 4.865000 2.635000 ;
      RECT 5.035000  0.255000 5.205000 0.615000 ;
      RECT 5.035000  2.105000 5.205000 2.465000 ;
      RECT 5.250000  0.955000 5.935000 1.125000 ;
      RECT 5.420000  0.765000 5.935000 0.955000 ;
      RECT 5.485000  2.125000 6.685000 2.465000 ;
      RECT 5.540000  0.255000 6.550000 0.505000 ;
      RECT 5.540000  0.505000 5.710000 0.595000 ;
      RECT 6.380000  0.505000 6.550000 0.655000 ;
      RECT 6.380000  0.655000 7.300000 0.825000 ;
      RECT 6.515000  1.935000 7.180000 2.105000 ;
      RECT 6.515000  2.105000 6.685000 2.125000 ;
      RECT 6.780000  0.085000 7.110000 0.445000 ;
      RECT 6.890000  2.275000 7.220000 2.635000 ;
      RECT 7.010000  1.470000 7.300000 1.640000 ;
      RECT 7.010000  1.640000 7.180000 1.935000 ;
      RECT 7.130000  0.825000 7.300000 1.075000 ;
      RECT 7.130000  1.075000 7.800000 1.245000 ;
      RECT 7.130000  1.245000 7.300000 1.470000 ;
      RECT 7.815000  1.795000 7.985000 2.635000 ;
      RECT 7.895000  0.085000 8.065000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  0.765000 2.155000 0.935000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 5.685000  0.765000 5.855000 0.935000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 1.925000 0.735000 2.215000 0.780000 ;
      RECT 1.925000 0.780000 5.915000 0.920000 ;
      RECT 1.925000 0.920000 2.215000 0.965000 ;
      RECT 5.625000 0.735000 5.915000 0.780000 ;
      RECT 5.625000 0.920000 5.915000 0.965000 ;
  END
END sky130_fd_sc_hd__fa_2
MACRO sky130_fd_sc_hd__fa_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fa_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 0.995000 1.240000 1.275000 ;
        RECT 0.910000 1.275000 1.080000 1.325000 ;
      LAYER mcon ;
        RECT 1.070000 1.105000 1.240000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.230000 1.030000 2.620000 1.360000 ;
      LAYER mcon ;
        RECT 2.450000 1.105000 2.620000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.250000 0.955000 4.625000 1.275000 ;
      LAYER mcon ;
        RECT 4.310000 1.105000 4.480000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.885000 1.035000 6.325000 1.275000 ;
      LAYER mcon ;
        RECT 6.150000 1.105000 6.320000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.010000 1.075000 1.300000 1.120000 ;
        RECT 1.010000 1.120000 6.380000 1.260000 ;
        RECT 1.010000 1.260000 1.300000 1.305000 ;
        RECT 2.390000 1.075000 2.680000 1.120000 ;
        RECT 2.390000 1.260000 2.680000 1.305000 ;
        RECT 4.250000 1.075000 4.540000 1.120000 ;
        RECT 4.250000 1.260000 4.540000 1.305000 ;
        RECT 6.090000 1.075000 6.380000 1.120000 ;
        RECT 6.090000 1.260000 6.380000 1.305000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.300000 1.445000 1.700000 1.880000 ;
      LAYER mcon ;
        RECT 1.530000 1.445000 1.700000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.200000 1.435000 3.560000 1.765000 ;
      LAYER mcon ;
        RECT 3.390000 1.445000 3.560000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.635000 1.445000 6.055000 1.765000 ;
      LAYER mcon ;
        RECT 5.690000 1.445000 5.860000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.470000 1.415000 1.760000 1.460000 ;
        RECT 1.470000 1.460000 5.920000 1.600000 ;
        RECT 1.470000 1.600000 1.760000 1.645000 ;
        RECT 3.330000 1.415000 3.620000 1.460000 ;
        RECT 3.330000 1.600000 3.620000 1.645000 ;
        RECT 5.630000 1.415000 5.920000 1.460000 ;
        RECT 5.630000 1.600000 5.920000 1.645000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.670000 1.105000 2.040000 1.275000 ;
        RECT 1.870000 1.275000 2.040000 1.595000 ;
        RECT 1.870000 1.595000 2.960000 1.765000 ;
        RECT 2.790000 0.965000 3.955000 1.250000 ;
        RECT 2.790000 1.250000 2.960000 1.595000 ;
        RECT 3.785000 1.250000 3.955000 1.515000 ;
        RECT 3.785000 1.515000 5.405000 1.685000 ;
        RECT 5.155000 1.685000 5.405000 1.955000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.345000 0.830000 ;
        RECT 0.085000 0.830000 0.260000 1.485000 ;
        RECT 0.085000 1.485000 0.345000 2.465000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.840000 0.255000 7.240000 0.810000 ;
        RECT 6.840000 1.485000 7.240000 2.465000 ;
        RECT 6.910000 0.810000 7.240000 1.485000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.430000  0.995000 0.685000 1.325000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  0.635000 1.710000 0.805000 ;
      RECT 0.515000  0.805000 0.685000 0.995000 ;
      RECT 0.515000  1.325000 0.685000 1.625000 ;
      RECT 0.515000  1.625000 1.105000 1.945000 ;
      RECT 0.515000  2.150000 0.765000 2.635000 ;
      RECT 0.935000  1.945000 1.105000 2.065000 ;
      RECT 0.935000  2.065000 1.710000 2.465000 ;
      RECT 1.110000  0.255000 1.710000 0.635000 ;
      RECT 1.470000  0.805000 1.710000 0.935000 ;
      RECT 1.960000  0.255000 2.130000 0.615000 ;
      RECT 1.960000  0.615000 2.970000 0.785000 ;
      RECT 1.960000  1.935000 3.035000 2.105000 ;
      RECT 1.960000  2.105000 2.130000 2.465000 ;
      RECT 2.300000  0.085000 2.630000 0.445000 ;
      RECT 2.300000  2.275000 2.630000 2.635000 ;
      RECT 2.800000  0.255000 2.970000 0.615000 ;
      RECT 2.800000  2.105000 3.035000 2.465000 ;
      RECT 3.240000  0.085000 3.570000 0.490000 ;
      RECT 3.240000  2.255000 3.570000 2.635000 ;
      RECT 3.740000  0.255000 3.910000 0.615000 ;
      RECT 3.740000  0.615000 4.750000 0.785000 ;
      RECT 3.740000  1.935000 4.750000 2.105000 ;
      RECT 3.740000  2.105000 3.910000 2.465000 ;
      RECT 4.080000  0.085000 4.410000 0.445000 ;
      RECT 4.080000  2.275000 4.410000 2.635000 ;
      RECT 4.580000  0.255000 4.750000 0.615000 ;
      RECT 4.580000  2.105000 4.750000 2.465000 ;
      RECT 4.795000  0.955000 5.460000 1.125000 ;
      RECT 4.965000  0.765000 5.460000 0.955000 ;
      RECT 5.085000  0.255000 6.095000 0.505000 ;
      RECT 5.085000  0.505000 5.255000 0.595000 ;
      RECT 5.085000  2.125000 6.170000 2.465000 ;
      RECT 5.925000  0.505000 6.095000 0.615000 ;
      RECT 5.925000  0.615000 6.665000 0.785000 ;
      RECT 6.000000  1.935000 6.665000 2.105000 ;
      RECT 6.000000  2.105000 6.170000 2.125000 ;
      RECT 6.265000  0.085000 6.595000 0.445000 ;
      RECT 6.340000  2.275000 6.670000 2.635000 ;
      RECT 6.495000  0.785000 6.665000 0.995000 ;
      RECT 6.495000  0.995000 6.740000 1.325000 ;
      RECT 6.495000  1.325000 6.665000 1.935000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.530000  0.765000 1.700000 0.935000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.230000  0.765000 5.400000 0.935000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
    LAYER met1 ;
      RECT 1.470000 0.735000 1.760000 0.780000 ;
      RECT 1.470000 0.780000 5.460000 0.920000 ;
      RECT 1.470000 0.920000 1.760000 0.965000 ;
      RECT 5.170000 0.735000 5.460000 0.780000 ;
      RECT 5.170000 0.920000 5.460000 0.965000 ;
  END
END sky130_fd_sc_hd__fa_1
MACRO sky130_fd_sc_hd__fa_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fa_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.633000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.080000 0.995000 2.680000 1.275000 ;
        RECT 2.080000 1.275000 2.340000 1.325000 ;
      LAYER mcon ;
        RECT 2.450000 1.105000 2.620000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.610000 1.030000 4.000000 1.360000 ;
      LAYER mcon ;
        RECT 3.830000 1.105000 4.000000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.645000 0.955000 6.005000 1.275000 ;
      LAYER mcon ;
        RECT 5.690000 1.105000 5.860000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.030000 0.995000 7.885000 1.275000 ;
      LAYER mcon ;
        RECT 7.070000 1.105000 7.240000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.390000 1.075000 2.680000 1.120000 ;
        RECT 2.390000 1.120000 7.300000 1.260000 ;
        RECT 2.390000 1.260000 2.680000 1.305000 ;
        RECT 3.770000 1.075000 4.060000 1.120000 ;
        RECT 3.770000 1.260000 4.060000 1.305000 ;
        RECT 5.630000 1.075000 5.920000 1.120000 ;
        RECT 5.630000 1.260000 5.920000 1.305000 ;
        RECT 7.010000 1.075000 7.300000 1.120000 ;
        RECT 7.010000 1.260000 7.300000 1.305000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.633000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.480000 1.445000 3.080000 1.690000 ;
      LAYER mcon ;
        RECT 2.910000 1.445000 3.080000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.580000 1.435000 4.995000 1.745000 ;
      LAYER mcon ;
        RECT 4.770000 1.445000 4.940000 1.615000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.075000 1.445000 7.760000 1.735000 ;
      LAYER mcon ;
        RECT 7.530000 1.445000 7.700000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.850000 1.415000 3.140000 1.460000 ;
        RECT 2.850000 1.460000 7.760000 1.600000 ;
        RECT 2.850000 1.600000 3.140000 1.645000 ;
        RECT 4.710000 1.415000 5.000000 1.460000 ;
        RECT 4.710000 1.600000 5.000000 1.645000 ;
        RECT 7.470000 1.415000 7.760000 1.460000 ;
        RECT 7.470000 1.600000 7.760000 1.645000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.477000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.050000 1.105000 3.420000 1.275000 ;
        RECT 3.250000 1.275000 3.420000 1.570000 ;
        RECT 3.250000 1.570000 4.340000 1.740000 ;
        RECT 4.170000 0.965000 5.390000 1.250000 ;
        RECT 4.170000 1.250000 4.340000 1.570000 ;
        RECT 5.220000 1.250000 5.390000 1.435000 ;
        RECT 5.220000 1.435000 5.580000 1.515000 ;
        RECT 5.220000 1.515000 6.845000 1.685000 ;
        RECT 6.595000 1.355000 6.845000 1.515000 ;
        RECT 6.595000 1.685000 6.845000 1.955000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.735000 1.525000 0.905000 ;
        RECT 0.085000 0.905000 0.435000 1.415000 ;
        RECT 0.085000 1.415000 1.570000 1.585000 ;
        RECT 0.515000 0.255000 0.845000 0.735000 ;
        RECT 0.515000 1.585000 0.845000 2.445000 ;
        RECT 1.355000 0.315000 1.685000 0.485000 ;
        RECT 1.355000 0.485000 1.525000 0.735000 ;
        RECT 1.400000 1.585000 1.570000 1.780000 ;
        RECT 1.400000 1.780000 1.645000 1.950000 ;
        RECT 1.435000 1.950000 1.645000 2.465000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.943000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.320000 0.255000  8.650000 0.485000 ;
        RECT 8.320000 1.795000  8.570000 1.965000 ;
        RECT 8.320000 1.965000  8.490000 2.465000 ;
        RECT 8.400000 0.485000  8.650000 0.735000 ;
        RECT 8.400000 0.735000 10.035000 0.905000 ;
        RECT 8.400000 1.415000 10.035000 1.585000 ;
        RECT 8.400000 1.585000  8.570000 1.795000 ;
        RECT 9.160000 0.270000  9.490000 0.735000 ;
        RECT 9.160000 1.585000  9.490000 2.425000 ;
        RECT 9.700000 0.905000 10.035000 1.415000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.175000  0.085000  0.345000 0.565000 ;
      RECT 0.175000  1.795000  0.345000 2.635000 ;
      RECT 0.605000  1.075000  1.910000 1.245000 ;
      RECT 1.015000  0.085000  1.185000 0.565000 ;
      RECT 1.015000  1.795000  1.185000 2.635000 ;
      RECT 1.740000  0.655000  3.090000 0.825000 ;
      RECT 1.740000  0.825000  1.910000 1.075000 ;
      RECT 1.740000  1.245000  1.910000 1.430000 ;
      RECT 1.740000  1.430000  1.945000 1.495000 ;
      RECT 1.740000  1.495000  2.310000 1.600000 ;
      RECT 1.775000  1.600000  2.310000 1.665000 ;
      RECT 1.815000  2.275000  2.145000 2.635000 ;
      RECT 1.855000  0.085000  2.185000 0.465000 ;
      RECT 2.140000  1.665000  2.310000 1.910000 ;
      RECT 2.140000  1.910000  3.170000 2.080000 ;
      RECT 2.370000  0.255000  3.090000 0.655000 ;
      RECT 2.735000  2.080000  3.170000 2.465000 ;
      RECT 2.850000  0.825000  3.090000 0.935000 ;
      RECT 3.340000  0.255000  3.510000 0.615000 ;
      RECT 3.340000  0.615000  4.350000 0.785000 ;
      RECT 3.340000  1.935000  4.415000 2.105000 ;
      RECT 3.340000  2.105000  3.510000 2.465000 ;
      RECT 3.680000  0.085000  4.010000 0.445000 ;
      RECT 3.680000  2.275000  4.010000 2.635000 ;
      RECT 4.180000  0.255000  4.350000 0.615000 ;
      RECT 4.180000  2.105000  4.415000 2.465000 ;
      RECT 4.620000  0.085000  4.950000 0.490000 ;
      RECT 4.620000  1.915000  4.950000 2.635000 ;
      RECT 5.120000  0.255000  5.290000 0.615000 ;
      RECT 5.120000  0.615000  6.130000 0.785000 ;
      RECT 5.120000  1.935000  6.130000 2.105000 ;
      RECT 5.120000  2.105000  5.290000 2.465000 ;
      RECT 5.460000  0.085000  5.790000 0.445000 ;
      RECT 5.460000  2.275000  5.790000 2.635000 ;
      RECT 5.960000  0.255000  6.130000 0.615000 ;
      RECT 5.960000  2.105000  6.130000 2.465000 ;
      RECT 6.175000  0.955000  6.860000 1.125000 ;
      RECT 6.345000  0.765000  6.860000 0.955000 ;
      RECT 6.410000  2.125000  7.610000 2.465000 ;
      RECT 6.465000  0.255000  7.475000 0.505000 ;
      RECT 6.465000  0.505000  6.635000 0.595000 ;
      RECT 7.305000  0.505000  7.475000 0.655000 ;
      RECT 7.305000  0.655000  8.225000 0.825000 ;
      RECT 7.440000  1.935000  8.105000 2.105000 ;
      RECT 7.440000  2.105000  7.610000 2.125000 ;
      RECT 7.705000  0.085000  8.035000 0.445000 ;
      RECT 7.815000  2.275000  8.145000 2.635000 ;
      RECT 7.935000  1.470000  8.225000 1.640000 ;
      RECT 7.935000  1.640000  8.105000 1.935000 ;
      RECT 8.055000  0.825000  8.225000 1.075000 ;
      RECT 8.055000  1.075000  9.445000 1.245000 ;
      RECT 8.055000  1.245000  8.225000 1.470000 ;
      RECT 8.740000  1.795000  8.910000 2.635000 ;
      RECT 8.820000  0.085000  8.990000 0.565000 ;
      RECT 9.660000  0.085000  9.830000 0.565000 ;
      RECT 9.660000  1.795000  9.830000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.910000  0.765000 3.080000 0.935000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 6.610000  0.765000 6.780000 0.935000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 2.850000 0.735000 3.140000 0.780000 ;
      RECT 2.850000 0.780000 6.840000 0.920000 ;
      RECT 2.850000 0.920000 3.140000 0.965000 ;
      RECT 6.550000 0.735000 6.840000 0.780000 ;
      RECT 6.550000 0.920000 6.840000 0.965000 ;
  END
END sky130_fd_sc_hd__fa_4
MACRO sky130_fd_sc_hd__clkdlybuf4s50_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s50_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.535000 1.290000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.190000 0.255000 3.595000 0.640000 ;
        RECT 3.190000 1.690000 3.595000 2.465000 ;
        RECT 3.345000 0.640000 3.595000 1.690000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.255000 0.415000 0.735000 ;
      RECT 0.085000  0.735000 1.055000 0.905000 ;
      RECT 0.085000  1.460000 1.055000 1.630000 ;
      RECT 0.085000  1.630000 0.430000 2.465000 ;
      RECT 0.585000  0.085000 0.915000 0.565000 ;
      RECT 0.600000  1.800000 0.930000 2.635000 ;
      RECT 0.705000  0.905000 1.055000 1.025000 ;
      RECT 0.705000  1.025000 1.135000 1.315000 ;
      RECT 0.705000  1.315000 1.055000 1.460000 ;
      RECT 1.380000  0.255000 1.730000 1.070000 ;
      RECT 1.380000  1.070000 2.240000 1.320000 ;
      RECT 1.380000  1.320000 1.730000 2.465000 ;
      RECT 1.990000  0.255000 2.240000 0.730000 ;
      RECT 1.990000  0.730000 2.580000 0.900000 ;
      RECT 1.990000  1.495000 2.580000 1.665000 ;
      RECT 1.990000  1.665000 2.240000 2.465000 ;
      RECT 2.410000  0.900000 2.580000 0.995000 ;
      RECT 2.410000  0.995000 3.175000 1.325000 ;
      RECT 2.410000  1.325000 2.580000 1.495000 ;
      RECT 2.690000  0.085000 3.020000 0.600000 ;
      RECT 2.690000  1.835000 3.020000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s50_1
MACRO sky130_fd_sc_hd__clkdlybuf4s50_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s50_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.480000 1.285000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.390500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.185000 0.270000 3.625000 0.640000 ;
        RECT 3.185000 1.530000 3.625000 2.465000 ;
        RECT 3.345000 0.640000 3.625000 1.530000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.270000 0.415000 0.735000 ;
      RECT 0.085000  0.735000 1.270000 0.905000 ;
      RECT 0.085000  1.455000 1.270000 1.630000 ;
      RECT 0.085000  1.630000 0.430000 2.465000 ;
      RECT 0.585000  0.085000 0.915000 0.565000 ;
      RECT 0.600000  1.800000 0.930000 2.635000 ;
      RECT 0.765000  1.075000 1.435000 1.245000 ;
      RECT 0.850000  0.905000 1.270000 1.075000 ;
      RECT 0.850000  1.245000 1.270000 1.455000 ;
      RECT 1.390000  1.785000 1.795000 2.465000 ;
      RECT 1.440000  0.270000 1.795000 0.900000 ;
      RECT 1.625000  0.900000 1.795000 1.075000 ;
      RECT 1.625000  1.075000 2.305000 1.245000 ;
      RECT 1.625000  1.245000 1.795000 1.785000 ;
      RECT 1.985000  0.270000 2.235000 0.735000 ;
      RECT 1.985000  0.735000 2.645000 0.905000 ;
      RECT 1.985000  1.460000 2.645000 1.630000 ;
      RECT 1.985000  1.630000 2.235000 2.465000 ;
      RECT 2.475000  0.905000 2.645000 0.995000 ;
      RECT 2.475000  0.995000 3.175000 1.325000 ;
      RECT 2.475000  1.325000 2.645000 1.460000 ;
      RECT 2.685000  0.085000 3.015000 0.565000 ;
      RECT 2.685000  1.800000 3.015000 2.635000 ;
      RECT 3.795000  0.085000 4.055000 0.635000 ;
      RECT 3.795000  1.800000 4.055000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s50_2
MACRO sky130_fd_sc_hd__xnor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.255000 1.075000 2.705000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485000 1.075000 0.960000 1.285000 ;
        RECT 0.790000 1.285000 0.960000 1.445000 ;
        RECT 0.790000 1.445000 3.100000 1.615000 ;
        RECT 2.930000 1.075000 3.955000 1.285000 ;
        RECT 2.930000 1.285000 3.100000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.913000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.795000 5.295000 1.965000 ;
        RECT 3.725000 1.965000 3.935000 2.125000 ;
        RECT 4.585000 0.305000 5.895000 0.475000 ;
        RECT 5.045000 1.415000 5.895000 1.625000 ;
        RECT 5.045000 1.625000 5.295000 1.795000 ;
        RECT 5.045000 1.965000 5.295000 2.125000 ;
        RECT 5.505000 0.475000 5.895000 1.415000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.085000  0.645000 0.860000 0.895000 ;
      RECT 0.085000  0.895000 0.315000 1.785000 ;
      RECT 0.085000  1.785000 3.480000 1.955000 ;
      RECT 0.085000  1.955000 2.080000 1.965000 ;
      RECT 0.085000  1.965000 0.400000 2.465000 ;
      RECT 0.105000  0.255000 1.280000 0.475000 ;
      RECT 0.570000  2.135000 0.820000 2.635000 ;
      RECT 0.990000  1.965000 1.240000 2.465000 ;
      RECT 1.030000  0.475000 1.280000 0.725000 ;
      RECT 1.030000  0.725000 2.120000 0.905000 ;
      RECT 1.410000  2.135000 1.660000 2.635000 ;
      RECT 1.450000  0.085000 1.620000 0.555000 ;
      RECT 1.790000  0.255000 2.120000 0.725000 ;
      RECT 1.830000  1.965000 2.080000 2.465000 ;
      RECT 2.390000  2.125000 2.640000 2.465000 ;
      RECT 2.430000  0.085000 2.600000 0.905000 ;
      RECT 2.770000  0.255000 3.100000 0.725000 ;
      RECT 2.770000  0.725000 5.335000 0.905000 ;
      RECT 2.810000  2.135000 3.060000 2.635000 ;
      RECT 3.230000  2.125000 3.555000 2.295000 ;
      RECT 3.230000  2.295000 4.355000 2.465000 ;
      RECT 3.270000  0.085000 3.440000 0.555000 ;
      RECT 3.310000  1.455000 4.805000 1.625000 ;
      RECT 3.310000  1.625000 3.480000 1.785000 ;
      RECT 3.610000  0.255000 3.975000 0.725000 ;
      RECT 4.105000  2.135000 4.355000 2.295000 ;
      RECT 4.145000  0.085000 4.315000 0.555000 ;
      RECT 4.625000  2.135000 4.875000 2.635000 ;
      RECT 4.635000  1.075000 5.295000 1.245000 ;
      RECT 4.635000  1.245000 4.805000 1.455000 ;
      RECT 5.005000  0.645000 5.335000 0.725000 ;
      RECT 5.465000  1.795000 5.895000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.465000  2.125000 2.635000 2.295000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.385000  2.125000 3.555000 2.295000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 2.405000 2.095000 2.695000 2.140000 ;
      RECT 2.405000 2.140000 3.615000 2.280000 ;
      RECT 2.405000 2.280000 2.695000 2.325000 ;
      RECT 3.325000 2.095000 3.615000 2.140000 ;
      RECT 3.325000 2.280000 3.615000 2.325000 ;
  END
END sky130_fd_sc_hd__xnor2_2
MACRO sky130_fd_sc_hd__xnor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.175000 1.075000 5.390000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 1.075000 1.855000 1.275000 ;
        RECT 1.685000 1.275000 1.855000 1.445000 ;
        RECT 1.685000 1.445000 5.730000 1.615000 ;
        RECT 5.560000 1.075000 7.430000 1.275000 ;
        RECT 5.560000 1.275000 5.730000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.721000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.160000 1.785000  8.250000 2.045000 ;
        RECT 7.960000 1.445000 10.035000 1.665000 ;
        RECT 7.960000 1.665000  8.250000 1.785000 ;
        RECT 7.960000 2.045000  8.250000 2.465000 ;
        RECT 8.380000 0.645000 10.035000 0.905000 ;
        RECT 8.840000 1.665000  9.090000 2.465000 ;
        RECT 9.680000 1.665000 10.035000 2.465000 ;
        RECT 9.815000 0.905000 10.035000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.645000  1.760000 0.905000 ;
      RECT 0.085000  0.905000  0.320000 1.445000 ;
      RECT 0.085000  1.445000  1.300000 1.615000 ;
      RECT 0.085000  1.615000  0.460000 2.465000 ;
      RECT 0.170000  0.255000  2.180000 0.475000 ;
      RECT 0.630000  1.835000  0.880000 2.635000 ;
      RECT 1.050000  1.615000  1.300000 1.785000 ;
      RECT 1.050000  1.785000  3.820000 2.005000 ;
      RECT 1.050000  2.005000  1.300000 2.465000 ;
      RECT 1.470000  2.175000  1.720000 2.635000 ;
      RECT 1.890000  2.005000  2.140000 2.465000 ;
      RECT 1.930000  0.475000  2.180000 0.725000 ;
      RECT 1.930000  0.725000  3.860000 0.905000 ;
      RECT 2.310000  2.175000  2.560000 2.635000 ;
      RECT 2.350000  0.085000  2.520000 0.555000 ;
      RECT 2.690000  0.255000  3.020000 0.725000 ;
      RECT 2.730000  2.005000  2.980000 2.465000 ;
      RECT 3.150000  2.175000  3.400000 2.635000 ;
      RECT 3.190000  0.085000  3.360000 0.555000 ;
      RECT 3.530000  0.255000  3.860000 0.725000 ;
      RECT 3.570000  2.005000  3.820000 2.465000 ;
      RECT 4.035000  0.085000  4.310000 0.905000 ;
      RECT 4.035000  1.785000  5.990000 2.005000 ;
      RECT 4.035000  2.005000  4.350000 2.465000 ;
      RECT 4.480000  0.255000  4.810000 0.725000 ;
      RECT 4.480000  0.725000  7.430000 0.735000 ;
      RECT 4.480000  0.735000  8.210000 0.905000 ;
      RECT 4.520000  2.175000  4.770000 2.635000 ;
      RECT 4.940000  2.005000  5.190000 2.465000 ;
      RECT 4.980000  0.085000  5.150000 0.555000 ;
      RECT 5.320000  0.255000  5.650000 0.725000 ;
      RECT 5.360000  2.175000  5.610000 2.635000 ;
      RECT 5.780000  2.005000  5.990000 2.215000 ;
      RECT 5.780000  2.215000  7.750000 2.465000 ;
      RECT 5.820000  0.085000  5.990000 0.555000 ;
      RECT 5.900000  1.445000  7.770000 1.615000 ;
      RECT 6.160000  0.255000  6.490000 0.725000 ;
      RECT 6.660000  0.085000  6.830000 0.555000 ;
      RECT 7.000000  0.255000  7.330000 0.725000 ;
      RECT 7.500000  0.085000  7.770000 0.555000 ;
      RECT 7.600000  1.075000  9.645000 1.275000 ;
      RECT 7.600000  1.275000  7.770000 1.445000 ;
      RECT 7.960000  0.305000  9.970000 0.475000 ;
      RECT 7.960000  0.475000  8.210000 0.735000 ;
      RECT 8.420000  1.835000  8.670000 2.635000 ;
      RECT 9.260000  1.835000  9.510000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  1.445000 1.235000 1.615000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  1.445000 6.295000 1.615000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
    LAYER met1 ;
      RECT 1.005000 1.415000 1.295000 1.460000 ;
      RECT 1.005000 1.460000 6.355000 1.600000 ;
      RECT 1.005000 1.600000 1.295000 1.645000 ;
      RECT 6.065000 1.415000 6.355000 1.460000 ;
      RECT 6.065000 1.600000 6.355000 1.645000 ;
  END
END sky130_fd_sc_hd__xnor2_4
MACRO sky130_fd_sc_hd__xnor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.930000 1.075000 1.625000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.670000 1.445000 ;
        RECT 0.425000 1.445000 1.965000 1.615000 ;
        RECT 1.795000 1.075000 2.395000 1.245000 ;
        RECT 1.795000 1.245000 1.965000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.525000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265000 2.125000 2.645000 2.295000 ;
        RECT 2.475000 1.755000 3.135000 1.955000 ;
        RECT 2.475000 1.955000 2.645000 2.125000 ;
        RECT 2.815000 0.345000 3.135000 0.825000 ;
        RECT 2.965000 0.825000 3.135000 1.755000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.280000 0.550000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.785000 ;
      RECT 0.085000  1.785000 2.305000 1.955000 ;
      RECT 0.085000  2.125000 0.385000 2.635000 ;
      RECT 0.555000  1.955000 0.885000 2.465000 ;
      RECT 1.055000  0.085000 1.225000 0.905000 ;
      RECT 1.055000  2.125000 1.685000 2.635000 ;
      RECT 1.395000  0.255000 1.725000 0.735000 ;
      RECT 1.395000  0.735000 2.645000 0.825000 ;
      RECT 1.395000  0.825000 2.305000 0.905000 ;
      RECT 1.895000  0.085000 2.245000 0.475000 ;
      RECT 2.135000  0.655000 2.645000 0.735000 ;
      RECT 2.135000  1.415000 2.795000 1.585000 ;
      RECT 2.135000  1.585000 2.305000 1.785000 ;
      RECT 2.415000  0.255000 2.645000 0.655000 ;
      RECT 2.625000  0.995000 2.795000 1.415000 ;
      RECT 2.815000  2.125000 3.115000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__xnor2_1
MACRO sky130_fd_sc_hd__dlymetal6s2s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s2s_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.570000 1.700000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245000 0.255000 1.670000 0.825000 ;
        RECT 1.245000 1.495000 2.150000 1.675000 ;
        RECT 1.245000 1.675000 1.670000 2.465000 ;
        RECT 1.320000 0.825000 1.670000 0.995000 ;
        RECT 1.320000 0.995000 2.150000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120000 -0.085000 0.290000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.255000 0.520000 0.655000 ;
      RECT 0.085000  0.655000 1.075000 0.825000 ;
      RECT 0.085000  1.870000 1.075000 2.040000 ;
      RECT 0.085000  2.040000 0.520000 2.465000 ;
      RECT 0.690000  0.085000 1.075000 0.485000 ;
      RECT 0.690000  2.210000 1.075000 2.635000 ;
      RECT 0.740000  0.825000 1.075000 0.995000 ;
      RECT 0.740000  0.995000 1.150000 1.325000 ;
      RECT 0.740000  1.325000 1.075000 1.870000 ;
      RECT 1.840000  1.845000 2.670000 2.040000 ;
      RECT 1.840000  2.040000 2.115000 2.465000 ;
      RECT 1.860000  0.255000 2.115000 0.655000 ;
      RECT 1.860000  0.655000 2.670000 0.825000 ;
      RECT 2.285000  0.085000 2.670000 0.485000 ;
      RECT 2.285000  2.210000 2.670000 2.635000 ;
      RECT 2.320000  0.825000 2.670000 0.995000 ;
      RECT 2.320000  0.995000 2.745000 1.325000 ;
      RECT 2.320000  1.325000 2.670000 1.845000 ;
      RECT 2.840000  0.255000 3.085000 0.825000 ;
      RECT 2.840000  1.495000 3.565000 1.675000 ;
      RECT 2.840000  1.675000 3.085000 2.465000 ;
      RECT 2.915000  0.825000 3.085000 0.995000 ;
      RECT 2.915000  0.995000 3.565000 1.495000 ;
      RECT 3.275000  0.255000 3.530000 0.655000 ;
      RECT 3.275000  0.655000 4.085000 0.825000 ;
      RECT 3.275000  1.845000 4.085000 2.040000 ;
      RECT 3.275000  2.040000 3.530000 2.465000 ;
      RECT 3.700000  0.085000 4.085000 0.485000 ;
      RECT 3.700000  2.210000 4.085000 2.635000 ;
      RECT 3.735000  0.825000 4.085000 0.995000 ;
      RECT 3.735000  0.995000 4.160000 1.325000 ;
      RECT 3.735000  1.325000 4.085000 1.845000 ;
      RECT 4.255000  0.255000 4.515000 0.825000 ;
      RECT 4.255000  1.495000 4.515000 2.465000 ;
      RECT 4.330000  0.825000 4.515000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__dlymetal6s2s_1
MACRO sky130_fd_sc_hd__edfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__edfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.225000 0.255000 11.555000 2.420000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.400000 1.065000 9.845000 1.410000 ;
        RECT 9.400000 1.410000 9.730000 2.465000 ;
        RECT 9.515000 0.255000 9.845000 1.065000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.845000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.355000  0.255000  1.785000 0.515000 ;
      RECT  1.355000  0.515000  1.525000 1.890000 ;
      RECT  1.355000  1.890000  1.785000 2.465000 ;
      RECT  2.235000  0.085000  2.565000 0.515000 ;
      RECT  2.235000  1.890000  2.565000 2.635000 ;
      RECT  2.495000  1.355000  3.085000 1.720000 ;
      RECT  2.755000  1.720000  3.085000 2.425000 ;
      RECT  2.780000  0.255000  3.005000 0.845000 ;
      RECT  2.780000  0.845000  3.635000 1.175000 ;
      RECT  2.780000  1.175000  3.085000 1.355000 ;
      RECT  3.185000  0.085000  3.515000 0.610000 ;
      RECT  3.265000  1.825000  3.460000 2.635000 ;
      RECT  3.805000  0.685000  3.975000 1.320000 ;
      RECT  3.805000  1.320000  4.175000 1.650000 ;
      RECT  4.125000  1.820000  4.515000 2.020000 ;
      RECT  4.125000  2.020000  4.455000 2.465000 ;
      RECT  4.145000  0.255000  4.415000 0.980000 ;
      RECT  4.145000  0.980000  4.515000 1.150000 ;
      RECT  4.345000  1.150000  4.515000 1.820000 ;
      RECT  4.795000  1.125000  4.980000 1.720000 ;
      RECT  4.815000  0.735000  5.320000 0.955000 ;
      RECT  4.915000  2.175000  5.955000 2.375000 ;
      RECT  5.005000  0.255000  5.680000 0.565000 ;
      RECT  5.150000  0.955000  5.320000 1.655000 ;
      RECT  5.150000  1.655000  5.615000 2.005000 ;
      RECT  5.510000  0.565000  5.680000 1.315000 ;
      RECT  5.510000  1.315000  6.360000 1.485000 ;
      RECT  5.785000  1.485000  6.360000 1.575000 ;
      RECT  5.785000  1.575000  5.955000 2.175000 ;
      RECT  5.870000  0.765000  6.935000 1.045000 ;
      RECT  5.870000  1.045000  7.445000 1.065000 ;
      RECT  5.870000  1.065000  6.070000 1.095000 ;
      RECT  5.945000  0.085000  6.340000 0.560000 ;
      RECT  6.125000  1.835000  6.360000 2.635000 ;
      RECT  6.190000  1.245000  6.360000 1.315000 ;
      RECT  6.530000  0.255000  6.935000 0.765000 ;
      RECT  6.530000  1.065000  7.445000 1.375000 ;
      RECT  6.530000  1.375000  6.860000 2.465000 ;
      RECT  7.070000  2.105000  7.360000 2.635000 ;
      RECT  7.165000  0.085000  7.440000 0.615000 ;
      RECT  7.790000  1.245000  7.980000 1.965000 ;
      RECT  7.925000  2.165000  8.890000 2.355000 ;
      RECT  8.005000  0.705000  8.470000 1.035000 ;
      RECT  8.025000  0.330000  8.890000 0.535000 ;
      RECT  8.150000  1.035000  8.470000 1.995000 ;
      RECT  8.640000  0.535000  8.890000 2.165000 ;
      RECT  9.060000  1.495000  9.230000 2.635000 ;
      RECT  9.095000  0.085000  9.345000 0.900000 ;
      RECT  9.900000  1.575000 10.130000 2.010000 ;
      RECT 10.015000  0.890000 10.640000 1.220000 ;
      RECT 10.300000  0.255000 10.640000 0.890000 ;
      RECT 10.300000  1.220000 10.640000 2.465000 ;
      RECT 10.810000  0.085000 11.055000 0.900000 ;
      RECT 10.810000  1.465000 11.055000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.635000  1.785000  0.805000 1.955000 ;
      RECT  1.015000  1.445000  1.185000 1.615000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.355000  0.425000  1.525000 0.595000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.805000  0.765000  3.975000 0.935000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.185000  0.425000  4.355000 0.595000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.800000  1.445000  4.970000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.210000  1.785000  5.380000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.800000  1.785000  7.970000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.220000  1.445000  8.390000 1.615000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.680000  1.785000  8.850000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT  9.930000  1.785000 10.100000 1.955000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.390000  0.765000 10.560000 0.935000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000  8.030000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000  8.450000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 10.620000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.740000 1.415000  5.030000 1.460000 ;
      RECT  4.740000 1.600000  5.030000 1.645000 ;
      RECT  5.150000 1.755000  5.440000 1.800000 ;
      RECT  5.150000 1.940000  5.440000 1.985000 ;
      RECT  7.740000 1.755000  8.030000 1.800000 ;
      RECT  7.740000 1.940000  8.030000 1.985000 ;
      RECT  8.160000 1.415000  8.450000 1.460000 ;
      RECT  8.160000 1.600000  8.450000 1.645000 ;
      RECT  8.620000 1.755000  8.910000 1.800000 ;
      RECT  8.620000 1.800000 10.160000 1.940000 ;
      RECT  8.620000 1.940000  8.910000 1.985000 ;
      RECT  9.870000 1.755000 10.160000 1.800000 ;
      RECT  9.870000 1.940000 10.160000 1.985000 ;
      RECT 10.330000 0.735000 10.620000 0.780000 ;
      RECT 10.330000 0.920000 10.620000 0.965000 ;
  END
END sky130_fd_sc_hd__edfxbp_1
MACRO sky130_fd_sc_hd__or4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615000 0.995000 3.270000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.480000 2.125000 3.120000 2.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.995000 1.235000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.780000 0.415000 4.055000 0.760000 ;
        RECT 3.780000 1.495000 4.055000 2.465000 ;
        RECT 3.885000 0.760000 4.055000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.450000 0.400000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.865000 ;
      RECT 0.085000  1.865000 1.915000 2.035000 ;
      RECT 0.085000  2.035000 0.345000 2.455000 ;
      RECT 0.515000  2.205000 0.845000 2.635000 ;
      RECT 0.655000  0.085000 0.825000 0.825000 ;
      RECT 0.990000  1.525000 1.575000 1.695000 ;
      RECT 1.075000  0.450000 1.245000 0.655000 ;
      RECT 1.075000  0.655000 1.575000 0.825000 ;
      RECT 1.405000  0.825000 1.575000 1.075000 ;
      RECT 1.405000  1.075000 1.830000 1.245000 ;
      RECT 1.405000  1.245000 1.575000 1.525000 ;
      RECT 1.470000  0.085000 1.845000 0.485000 ;
      RECT 1.510000  2.205000 2.255000 2.375000 ;
      RECT 1.745000  1.415000 2.395000 1.585000 ;
      RECT 1.745000  1.585000 1.915000 1.865000 ;
      RECT 2.015000  0.305000 2.185000 0.655000 ;
      RECT 2.015000  0.655000 3.610000 0.825000 ;
      RECT 2.085000  1.785000 3.120000 1.955000 ;
      RECT 2.085000  1.955000 2.255000 2.205000 ;
      RECT 2.225000  0.995000 2.395000 1.415000 ;
      RECT 2.370000  0.085000 2.700000 0.485000 ;
      RECT 2.870000  0.305000 3.040000 0.655000 ;
      RECT 2.950000  1.495000 3.610000 1.665000 ;
      RECT 2.950000  1.665000 3.120000 1.785000 ;
      RECT 3.210000  0.085000 3.590000 0.485000 ;
      RECT 3.290000  1.835000 3.570000 2.635000 ;
      RECT 3.440000  0.825000 3.610000 0.995000 ;
      RECT 3.440000  0.995000 3.715000 1.325000 ;
      RECT 3.440000  1.325000 3.610000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__or4bb_1
MACRO sky130_fd_sc_hd__or4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.640000 0.995000 3.295000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 2.125000 3.145000 2.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.780000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.995000 1.240000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.415000 4.080000 0.760000 ;
        RECT 3.805000 1.495000 4.080000 2.465000 ;
        RECT 3.910000 0.760000 4.080000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.450000 0.405000 0.825000 ;
      RECT 0.085000  0.825000 0.260000 1.865000 ;
      RECT 0.085000  1.865000 1.940000 2.035000 ;
      RECT 0.085000  2.035000 0.345000 2.455000 ;
      RECT 0.515000  2.205000 0.845000 2.635000 ;
      RECT 0.660000  0.085000 0.830000 0.825000 ;
      RECT 0.995000  1.525000 1.600000 1.695000 ;
      RECT 1.080000  0.450000 1.250000 0.655000 ;
      RECT 1.080000  0.655000 1.600000 0.825000 ;
      RECT 1.410000  0.825000 1.600000 1.075000 ;
      RECT 1.410000  1.075000 1.855000 1.245000 ;
      RECT 1.410000  1.245000 1.600000 1.525000 ;
      RECT 1.495000  0.085000 1.850000 0.485000 ;
      RECT 1.535000  2.205000 2.280000 2.375000 ;
      RECT 1.770000  1.415000 2.420000 1.585000 ;
      RECT 1.770000  1.585000 1.940000 1.865000 ;
      RECT 2.025000  0.305000 2.195000 0.655000 ;
      RECT 2.025000  0.655000 3.635000 0.825000 ;
      RECT 2.110000  1.785000 3.145000 1.955000 ;
      RECT 2.110000  1.955000 2.280000 2.205000 ;
      RECT 2.250000  0.995000 2.420000 1.415000 ;
      RECT 2.395000  0.085000 2.725000 0.485000 ;
      RECT 2.895000  0.305000 3.065000 0.655000 ;
      RECT 2.975000  1.495000 3.635000 1.665000 ;
      RECT 2.975000  1.665000 3.145000 1.785000 ;
      RECT 3.235000  0.085000 3.615000 0.485000 ;
      RECT 3.315000  1.835000 3.595000 2.635000 ;
      RECT 3.465000  0.825000 3.635000 0.995000 ;
      RECT 3.465000  0.995000 3.740000 1.325000 ;
      RECT 3.465000  1.325000 3.635000 1.495000 ;
      RECT 4.250000  0.085000 4.420000 1.025000 ;
      RECT 4.250000  1.440000 4.420000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__or4bb_2
MACRO sky130_fd_sc_hd__or4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.235000 0.995000 3.405000 1.445000 ;
        RECT 3.235000 1.445000 3.670000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675000 0.995000 3.005000 1.450000 ;
        RECT 2.795000 1.450000 3.005000 1.785000 ;
        RECT 2.795000 1.785000 3.115000 2.375000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.695000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.995000 1.235000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.875000 1.455000 5.435000 1.625000 ;
        RECT 3.875000 1.625000 4.125000 2.465000 ;
        RECT 3.915000 0.255000 4.165000 0.725000 ;
        RECT 3.915000 0.725000 5.435000 0.905000 ;
        RECT 4.675000 0.255000 5.005000 0.725000 ;
        RECT 4.715000 1.625000 4.965000 2.465000 ;
        RECT 5.205000 0.905000 5.435000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.085000  0.450000 0.400000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.865000 ;
      RECT 0.085000  1.865000 1.295000 2.035000 ;
      RECT 0.085000  2.035000 0.345000 2.455000 ;
      RECT 0.515000  2.205000 0.845000 2.635000 ;
      RECT 0.655000  0.085000 0.825000 0.825000 ;
      RECT 0.990000  1.525000 1.595000 1.695000 ;
      RECT 1.075000  0.450000 1.245000 0.655000 ;
      RECT 1.075000  0.655000 1.595000 0.825000 ;
      RECT 1.125000  2.035000 1.295000 2.295000 ;
      RECT 1.125000  2.295000 2.445000 2.465000 ;
      RECT 1.405000  0.825000 1.595000 0.995000 ;
      RECT 1.405000  0.995000 1.695000 1.325000 ;
      RECT 1.405000  1.325000 1.595000 1.525000 ;
      RECT 1.510000  1.955000 2.105000 2.125000 ;
      RECT 1.515000  0.085000 1.845000 0.480000 ;
      RECT 1.935000  0.655000 3.745000 0.825000 ;
      RECT 1.935000  0.825000 2.105000 1.955000 ;
      RECT 2.095000  0.305000 2.265000 0.655000 ;
      RECT 2.275000  0.995000 2.445000 2.295000 ;
      RECT 2.465000  0.085000 2.795000 0.485000 ;
      RECT 2.965000  0.305000 3.135000 0.655000 ;
      RECT 3.355000  0.085000 3.735000 0.485000 ;
      RECT 3.400000  1.795000 3.650000 2.635000 ;
      RECT 3.575000  0.825000 3.745000 1.075000 ;
      RECT 3.575000  1.075000 5.035000 1.245000 ;
      RECT 4.295000  1.795000 4.545000 2.635000 ;
      RECT 4.335000  0.085000 4.505000 0.555000 ;
      RECT 5.135000  1.795000 5.385000 2.635000 ;
      RECT 5.175000  0.085000 5.345000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__or4bb_4
MACRO sky130_fd_sc_hd__tapvpwrvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvpwrvgnd_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
      LAYER pwell ;
        RECT 0.145000 0.320000 0.315000 0.845000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
      LAYER nwell ;
        RECT -0.190000 1.305000 0.650000 2.910000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.460000 0.085000 ;
      RECT 0.000000  2.635000 0.460000 2.805000 ;
      RECT 0.085000  0.085000 0.375000 0.810000 ;
      RECT 0.085000  1.470000 0.375000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
  END
END sky130_fd_sc_hd__tapvpwrvgnd_1
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.265000 1.065000 ;
        RECT 0.085000 1.065000 0.575000 1.285000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.270000 1.075000 8.010000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  2.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 0.255000 2.335000 0.725000 ;
        RECT 2.005000 0.725000 8.655000 0.905000 ;
        RECT 2.845000 0.255000 3.175000 0.725000 ;
        RECT 3.685000 0.255000 4.015000 0.725000 ;
        RECT 4.525000 0.255000 4.855000 0.725000 ;
        RECT 5.365000 0.255000 5.695000 0.725000 ;
        RECT 5.405000 1.445000 8.655000 1.615000 ;
        RECT 5.405000 1.615000 5.655000 2.125000 ;
        RECT 6.205000 0.255000 6.535000 0.725000 ;
        RECT 6.245000 1.615000 6.495000 2.125000 ;
        RECT 7.045000 0.255000 7.375000 0.725000 ;
        RECT 7.085000 1.615000 7.335000 2.125000 ;
        RECT 7.885000 0.255000 8.215000 0.725000 ;
        RECT 7.925000 1.615000 8.175000 2.125000 ;
        RECT 8.180000 0.905000 8.655000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.930000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.195000  1.455000 0.415000 2.635000 ;
      RECT 0.435000  0.085000 0.655000 0.895000 ;
      RECT 0.585000  1.455000 0.915000 2.465000 ;
      RECT 0.745000  1.065000 1.155000 1.075000 ;
      RECT 0.745000  1.075000 5.000000 1.285000 ;
      RECT 0.745000  1.285000 0.915000 1.455000 ;
      RECT 0.825000  0.255000 1.155000 1.065000 ;
      RECT 1.085000  1.455000 1.330000 2.635000 ;
      RECT 1.325000  0.085000 1.835000 0.905000 ;
      RECT 1.555000  1.455000 5.235000 1.665000 ;
      RECT 1.555000  1.665000 1.875000 2.465000 ;
      RECT 2.045000  1.835000 2.295000 2.635000 ;
      RECT 2.465000  1.665000 2.715000 2.465000 ;
      RECT 2.505000  0.085000 2.675000 0.555000 ;
      RECT 2.885000  1.835000 3.135000 2.635000 ;
      RECT 3.305000  1.665000 3.555000 2.465000 ;
      RECT 3.345000  0.085000 3.515000 0.555000 ;
      RECT 3.725000  1.835000 3.975000 2.635000 ;
      RECT 4.145000  1.665000 4.395000 2.465000 ;
      RECT 4.185000  0.085000 4.355000 0.555000 ;
      RECT 4.565000  1.835000 4.815000 2.635000 ;
      RECT 4.985000  1.665000 5.235000 2.295000 ;
      RECT 4.985000  2.295000 8.595000 2.465000 ;
      RECT 5.025000  0.085000 5.195000 0.555000 ;
      RECT 5.825000  1.785000 6.075000 2.295000 ;
      RECT 5.865000  0.085000 6.035000 0.555000 ;
      RECT 6.665000  1.785000 6.915000 2.295000 ;
      RECT 6.705000  0.085000 6.875000 0.555000 ;
      RECT 7.505000  1.785000 7.755000 2.295000 ;
      RECT 7.545000  0.085000 7.715000 0.555000 ;
      RECT 8.345000  1.785000 8.595000 2.295000 ;
      RECT 8.385000  0.085000 8.655000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_8
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.725000 0.325000 1.325000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 1.065000 1.325000 1.325000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.235000 0.255000 1.565000 0.725000 ;
        RECT 1.235000 0.725000 2.215000 0.895000 ;
        RECT 1.655000 1.850000 2.215000 2.465000 ;
        RECT 2.035000 0.895000 2.215000 1.850000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.330000  0.370000 0.675000 0.545000 ;
      RECT 0.415000  1.510000 1.705000 1.680000 ;
      RECT 0.415000  1.680000 0.675000 1.905000 ;
      RECT 0.495000  0.545000 0.675000 1.510000 ;
      RECT 0.855000  0.085000 1.065000 0.895000 ;
      RECT 0.875000  1.855000 1.205000 2.635000 ;
      RECT 1.535000  1.075000 1.865000 1.245000 ;
      RECT 1.535000  1.245000 1.705000 1.510000 ;
      RECT 1.735000  0.085000 2.120000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_1
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.56000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.315000 0.995000 ;
        RECT 0.085000 0.995000 0.665000 1.325000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  3.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.450000 1.075000 15.650000 1.285000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  4.968000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  2.925000 0.255000  3.255000 0.725000 ;
        RECT  2.925000 0.725000 16.475000 0.905000 ;
        RECT  3.765000 0.255000  4.095000 0.725000 ;
        RECT  4.605000 0.255000  4.935000 0.725000 ;
        RECT  5.445000 0.255000  5.775000 0.725000 ;
        RECT  6.285000 0.255000  6.615000 0.725000 ;
        RECT  7.125000 0.255000  7.455000 0.725000 ;
        RECT  7.965000 0.255000  8.295000 0.725000 ;
        RECT  8.805000 0.255000  9.135000 0.725000 ;
        RECT  9.645000 0.255000  9.975000 0.725000 ;
        RECT  9.685000 1.455000 16.475000 1.625000 ;
        RECT  9.685000 1.625000  9.935000 2.125000 ;
        RECT 10.485000 0.255000 10.815000 0.725000 ;
        RECT 10.525000 1.625000 10.775000 2.125000 ;
        RECT 11.325000 0.255000 11.655000 0.725000 ;
        RECT 11.365000 1.625000 11.615000 2.125000 ;
        RECT 12.165000 0.255000 12.495000 0.725000 ;
        RECT 12.205000 1.625000 12.455000 2.125000 ;
        RECT 13.005000 0.255000 13.335000 0.725000 ;
        RECT 13.045000 1.625000 13.295000 2.125000 ;
        RECT 13.845000 0.255000 14.175000 0.725000 ;
        RECT 13.885000 1.625000 14.135000 2.125000 ;
        RECT 14.685000 0.255000 15.015000 0.725000 ;
        RECT 14.725000 1.625000 14.975000 2.125000 ;
        RECT 15.525000 0.255000 15.855000 0.725000 ;
        RECT 15.565000 1.625000 15.815000 2.125000 ;
        RECT 15.820000 0.905000 16.475000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 16.560000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 16.750000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 16.560000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.560000 0.085000 ;
      RECT  0.000000  2.635000 16.560000 2.805000 ;
      RECT  0.300000  1.495000  0.515000 2.635000 ;
      RECT  0.485000  0.085000  0.815000 0.825000 ;
      RECT  0.685000  1.495000  1.015000 2.465000 ;
      RECT  0.835000  1.065000  2.035000 1.075000 ;
      RECT  0.835000  1.075000  9.280000 1.285000 ;
      RECT  0.835000  1.285000  1.015000 1.495000 ;
      RECT  0.985000  0.255000  1.195000 1.065000 ;
      RECT  1.185000  1.455000  1.355000 2.635000 ;
      RECT  1.365000  0.085000  1.615000 0.895000 ;
      RECT  1.525000  1.285000  1.855000 2.465000 ;
      RECT  1.785000  0.255000  2.035000 1.065000 ;
      RECT  2.025000  1.455000  2.270000 2.635000 ;
      RECT  2.205000  0.085000  2.755000 0.905000 ;
      RECT  2.475000  1.455000  9.515000 1.665000 ;
      RECT  2.475000  1.665000  2.795000 2.465000 ;
      RECT  2.965000  1.835000  3.215000 2.635000 ;
      RECT  3.385000  1.665000  3.635000 2.465000 ;
      RECT  3.425000  0.085000  3.595000 0.555000 ;
      RECT  3.805000  1.835000  4.055000 2.635000 ;
      RECT  4.225000  1.665000  4.475000 2.465000 ;
      RECT  4.265000  0.085000  4.435000 0.555000 ;
      RECT  4.645000  1.835000  4.895000 2.635000 ;
      RECT  5.065000  1.665000  5.315000 2.465000 ;
      RECT  5.105000  0.085000  5.275000 0.555000 ;
      RECT  5.485000  1.835000  5.735000 2.635000 ;
      RECT  5.905000  1.665000  6.155000 2.465000 ;
      RECT  5.945000  0.085000  6.115000 0.555000 ;
      RECT  6.325000  1.835000  6.575000 2.635000 ;
      RECT  6.745000  1.665000  6.995000 2.465000 ;
      RECT  6.785000  0.085000  6.955000 0.555000 ;
      RECT  7.165000  1.835000  7.415000 2.635000 ;
      RECT  7.585000  1.665000  7.835000 2.465000 ;
      RECT  7.625000  0.085000  7.795000 0.555000 ;
      RECT  8.005000  1.835000  8.255000 2.635000 ;
      RECT  8.425000  1.665000  8.675000 2.465000 ;
      RECT  8.465000  0.085000  8.635000 0.555000 ;
      RECT  8.845000  1.835000  9.095000 2.635000 ;
      RECT  9.265000  1.665000  9.515000 2.295000 ;
      RECT  9.265000  2.295000 16.235000 2.465000 ;
      RECT  9.305000  0.085000  9.475000 0.555000 ;
      RECT 10.105000  1.795000 10.355000 2.295000 ;
      RECT 10.145000  0.085000 10.315000 0.555000 ;
      RECT 10.945000  1.795000 11.195000 2.295000 ;
      RECT 10.985000  0.085000 11.155000 0.555000 ;
      RECT 11.785000  1.795000 12.035000 2.295000 ;
      RECT 11.825000  0.085000 11.995000 0.555000 ;
      RECT 12.625000  1.795000 12.875000 2.295000 ;
      RECT 12.665000  0.085000 12.835000 0.555000 ;
      RECT 13.465000  1.795000 13.715000 2.295000 ;
      RECT 13.505000  0.085000 13.675000 0.555000 ;
      RECT 14.305000  1.795000 14.555000 2.295000 ;
      RECT 14.345000  0.085000 14.515000 0.555000 ;
      RECT 15.145000  1.795000 15.395000 2.295000 ;
      RECT 15.185000  0.085000 15.355000 0.555000 ;
      RECT 15.985000  1.795000 16.235000 2.295000 ;
      RECT 16.025000  0.085000 16.295000 0.555000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_16
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.600000 1.065000 3.125000 1.275000 ;
        RECT 2.910000 1.275000 3.125000 1.965000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.480000 1.065000 0.920000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 1.705000 0.895000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 1.415000 0.895000 1.665000 2.125000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.895000 ;
      RECT 0.085000  1.445000 1.245000 1.655000 ;
      RECT 0.085000  1.655000 0.405000 2.465000 ;
      RECT 0.575000  1.825000 0.825000 2.635000 ;
      RECT 0.995000  1.655000 1.245000 2.295000 ;
      RECT 0.995000  2.295000 2.125000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.835000  1.445000 2.090000 1.890000 ;
      RECT 1.835000  1.890000 2.125000 2.295000 ;
      RECT 1.875000  0.085000 2.045000 0.895000 ;
      RECT 1.875000  1.075000 2.430000 1.245000 ;
      RECT 2.215000  0.725000 2.565000 0.895000 ;
      RECT 2.215000  0.895000 2.430000 1.075000 ;
      RECT 2.260000  1.245000 2.430000 1.445000 ;
      RECT 2.260000  1.445000 2.565000 1.615000 ;
      RECT 2.395000  0.445000 2.565000 0.725000 ;
      RECT 2.395000  1.615000 2.565000 2.460000 ;
      RECT 2.775000  0.085000 3.030000 0.845000 ;
      RECT 2.775000  2.145000 3.025000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_2
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.075000 4.975000 1.320000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.075000 1.800000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 3.385000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 2.295000 0.905000 2.625000 1.445000 ;
        RECT 2.295000 1.445000 3.305000 1.745000 ;
        RECT 2.295000 1.745000 2.465000 2.125000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 3.135000 1.745000 3.305000 2.125000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.085000 0.365000 0.905000 ;
      RECT 0.085000  1.455000 2.125000 1.665000 ;
      RECT 0.085000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.865000 2.635000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.035000  1.665000 1.205000 2.465000 ;
      RECT 1.375000  1.835000 1.625000 2.635000 ;
      RECT 1.795000  1.665000 2.125000 2.295000 ;
      RECT 1.795000  2.295000 3.855000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.635000  1.935000 2.965000 2.295000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 2.795000  1.075000 4.275000 1.275000 ;
      RECT 3.475000  1.575000 3.855000 2.295000 ;
      RECT 3.555000  0.085000 3.845000 0.905000 ;
      RECT 4.025000  0.255000 4.355000 0.815000 ;
      RECT 4.025000  0.815000 4.275000 1.075000 ;
      RECT 4.025000  1.275000 4.275000 1.575000 ;
      RECT 4.025000  1.575000 4.355000 2.465000 ;
      RECT 4.525000  0.085000 4.815000 0.905000 ;
      RECT 4.525000  1.495000 4.930000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_4
MACRO sky130_fd_sc_hd__a31oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 0.995000 2.665000 1.615000 ;
        RECT 2.905000 0.995000 3.075000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.995000 1.755000 1.615000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.995000 0.820000 1.615000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.820000 1.075000 4.490000 1.275000 ;
        RECT 4.265000 1.275000 4.490000 1.625000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.922000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 0.655000 4.505000 0.825000 ;
        RECT 3.255000 0.255000 3.425000 0.655000 ;
        RECT 3.255000 0.825000 3.570000 1.445000 ;
        RECT 3.255000 1.445000 4.085000 1.615000 ;
        RECT 3.755000 1.615000 4.085000 2.115000 ;
        RECT 4.175000 0.295000 4.505000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.095000  0.655000 2.105000 0.825000 ;
      RECT 0.175000  1.785000 3.505000 1.955000 ;
      RECT 0.175000  1.955000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.125000 0.845000 2.635000 ;
      RECT 1.015000  1.955000 1.185000 2.465000 ;
      RECT 1.355000  0.295000 3.075000 0.465000 ;
      RECT 1.355000  2.125000 1.685000 2.635000 ;
      RECT 1.855000  1.955000 2.025000 2.465000 ;
      RECT 2.310000  2.125000 2.980000 2.635000 ;
      RECT 3.335000  1.955000 3.505000 2.295000 ;
      RECT 3.335000  2.295000 4.425000 2.465000 ;
      RECT 3.675000  0.085000 4.005000 0.465000 ;
      RECT 4.255000  1.795000 4.425000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__a31oi_2
MACRO sky130_fd_sc_hd__a31oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 0.995000 5.420000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.995000 3.550000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.995000 1.735000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.670000 0.995000 6.855000 1.630000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.443500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.975000 0.635000 7.585000 0.805000 ;
        RECT 6.075000 1.915000 7.245000 2.085000 ;
        RECT 6.575000 0.255000 6.745000 0.635000 ;
        RECT 7.045000 0.805000 7.245000 1.915000 ;
        RECT 7.415000 0.255000 7.585000 0.635000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 3.785000 0.805000 ;
      RECT 0.175000  1.495000 5.405000 1.665000 ;
      RECT 0.175000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  1.915000 0.845000 2.635000 ;
      RECT 1.015000  0.255000 1.185000 0.635000 ;
      RECT 1.015000  1.665000 1.185000 2.465000 ;
      RECT 1.355000  0.085000 1.685000 0.465000 ;
      RECT 1.355000  1.915000 1.685000 2.635000 ;
      RECT 1.855000  0.255000 2.025000 0.635000 ;
      RECT 1.855000  1.665000 2.025000 2.465000 ;
      RECT 2.195000  0.295000 5.565000 0.465000 ;
      RECT 2.195000  1.915000 2.525000 2.635000 ;
      RECT 2.695000  1.665000 2.865000 2.465000 ;
      RECT 3.035000  1.915000 3.365000 2.635000 ;
      RECT 3.535000  1.665000 3.705000 2.465000 ;
      RECT 3.895000  1.915000 4.225000 2.635000 ;
      RECT 4.395000  1.665000 4.565000 2.465000 ;
      RECT 4.735000  2.255000 5.065000 2.635000 ;
      RECT 5.235000  1.665000 5.405000 2.255000 ;
      RECT 5.235000  2.255000 7.665000 2.425000 ;
      RECT 5.235000  2.425000 5.405000 2.465000 ;
      RECT 6.075000  0.085000 6.405000 0.465000 ;
      RECT 6.915000  0.085000 7.245000 0.465000 ;
      RECT 7.415000  1.495000 7.665000 2.255000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__a31oi_4
MACRO sky130_fd_sc_hd__a31oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.445000 1.455000 1.665000 ;
        RECT 1.270000 0.995000 1.455000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 0.335000 1.055000 1.275000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.365000 1.325000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 0.995000 2.215000 1.325000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.481250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.380000 0.295000 1.785000 0.715000 ;
        RECT 1.380000 0.715000 1.795000 0.825000 ;
        RECT 1.625000 0.825000 1.795000 1.495000 ;
        RECT 1.625000 1.495000 2.210000 1.665000 ;
        RECT 1.875000 1.665000 2.210000 2.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.090000  0.085000 0.430000 0.815000 ;
      RECT 0.090000  1.495000 0.420000 2.635000 ;
      RECT 0.590000  1.835000 1.695000 2.005000 ;
      RECT 0.590000  2.005000 0.765000 2.415000 ;
      RECT 0.935000  2.175000 1.265000 2.635000 ;
      RECT 1.470000  2.005000 1.695000 2.415000 ;
      RECT 1.955000  0.085000 2.215000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__a31oi_1
MACRO sky130_fd_sc_hd__a21boi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.545000 1.065000 4.970000 1.310000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.030000 1.065000 3.375000 1.480000 ;
        RECT 3.030000 1.480000 6.450000 1.705000 ;
        RECT 5.205000 1.075000 6.450000 1.480000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.075000 0.650000 1.615000 ;
        RECT 0.480000 0.995000 0.650000 1.075000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.288000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275000 0.370000 1.465000 0.615000 ;
        RECT 1.275000 0.615000 2.325000 0.695000 ;
        RECT 1.275000 0.695000 4.885000 0.865000 ;
        RECT 1.560000 1.585000 2.860000 1.705000 ;
        RECT 1.560000 1.705000 2.725000 2.035000 ;
        RECT 2.135000 0.255000 2.325000 0.615000 ;
        RECT 2.570000 0.865000 4.885000 0.895000 ;
        RECT 2.570000 0.895000 2.860000 1.585000 ;
        RECT 3.255000 0.675000 4.885000 0.695000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.090000  0.255000 0.445000 0.615000 ;
      RECT 0.090000  0.615000 1.105000 0.795000 ;
      RECT 0.125000  1.785000 0.990000 2.005000 ;
      RECT 0.125000  2.005000 0.455000 2.465000 ;
      RECT 0.625000  2.175000 0.885000 2.635000 ;
      RECT 0.720000  0.085000 1.105000 0.445000 ;
      RECT 0.820000  0.795000 1.105000 1.035000 ;
      RECT 0.820000  1.035000 2.400000 1.345000 ;
      RECT 0.820000  1.345000 0.990000 1.785000 ;
      RECT 1.160000  1.795000 1.355000 2.215000 ;
      RECT 1.160000  2.215000 3.095000 2.465000 ;
      RECT 1.635000  0.085000 1.965000 0.445000 ;
      RECT 1.935000  2.205000 3.095000 2.215000 ;
      RECT 2.495000  0.085000 3.085000 0.525000 ;
      RECT 2.895000  1.875000 6.605000 2.105000 ;
      RECT 2.895000  2.105000 3.095000 2.205000 ;
      RECT 3.265000  0.255000 5.315000 0.505000 ;
      RECT 3.265000  2.275000 3.595000 2.635000 ;
      RECT 4.125000  2.275000 4.455000 2.635000 ;
      RECT 4.625000  2.105000 4.815000 2.465000 ;
      RECT 4.985000  2.275000 5.315000 2.635000 ;
      RECT 5.055000  0.505000 5.315000 0.735000 ;
      RECT 5.055000  0.735000 6.175000 0.905000 ;
      RECT 5.485000  0.085000 5.675000 0.565000 ;
      RECT 5.485000  2.105000 5.665000 2.465000 ;
      RECT 5.845000  0.255000 6.175000 0.735000 ;
      RECT 5.845000  2.275000 6.175000 2.635000 ;
      RECT 6.345000  0.085000 6.605000 0.885000 ;
      RECT 6.345000  2.105000 6.605000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
END sky130_fd_sc_hd__a21boi_4
MACRO sky130_fd_sc_hd__a21boi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.605000 0.995000 3.215000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095000 1.075000 2.425000 1.245000 ;
        RECT 2.100000 1.245000 2.425000 1.495000 ;
        RECT 2.100000 1.495000 3.675000 1.675000 ;
        RECT 3.385000 1.035000 3.795000 1.295000 ;
        RECT 3.385000 1.295000 3.675000 1.495000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.765000 0.425000 1.805000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.627500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 0.255000 1.720000 0.615000 ;
        RECT 1.520000 0.615000 3.060000 0.785000 ;
        RECT 1.520000 0.785000 1.715000 2.115000 ;
        RECT 2.730000 0.255000 3.060000 0.615000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.095000  2.080000 0.425000 2.635000 ;
      RECT 0.265000  0.360000 0.795000 0.530000 ;
      RECT 0.595000  0.530000 0.795000 1.070000 ;
      RECT 0.595000  1.070000 1.325000 1.285000 ;
      RECT 0.595000  1.285000 0.855000 2.265000 ;
      RECT 0.985000  0.085000 1.225000 0.885000 ;
      RECT 1.045000  1.795000 1.350000 2.285000 ;
      RECT 1.045000  2.285000 2.215000 2.465000 ;
      RECT 1.885000  1.855000 3.920000 2.025000 ;
      RECT 1.885000  2.025000 2.215000 2.285000 ;
      RECT 1.940000  0.085000 2.270000 0.445000 ;
      RECT 2.385000  2.195000 2.555000 2.635000 ;
      RECT 2.810000  2.025000 3.920000 2.105000 ;
      RECT 2.810000  2.105000 2.980000 2.465000 ;
      RECT 3.160000  2.275000 3.490000 2.635000 ;
      RECT 3.635000  0.085000 3.930000 0.865000 ;
      RECT 3.660000  2.105000 3.920000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a21boi_2
MACRO sky130_fd_sc_hd__a21boi_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.765000 2.170000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.340000 0.765000 2.615000 1.435000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.470000 1.200000 0.895000 1.955000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.392200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.200000 1.610000 1.655000 ;
        RECT 1.065000 1.655000 1.305000 2.465000 ;
        RECT 1.315000 0.255000 1.610000 1.200000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  0.280000 0.380000 0.780000 ;
      RECT 0.095000  0.780000 1.145000 1.030000 ;
      RECT 0.095000  1.030000 0.300000 2.085000 ;
      RECT 0.095000  2.085000 0.355000 2.465000 ;
      RECT 0.525000  2.175000 0.855000 2.635000 ;
      RECT 0.550000  0.085000 1.145000 0.610000 ;
      RECT 1.475000  1.825000 2.665000 2.005000 ;
      RECT 1.475000  2.005000 1.805000 2.465000 ;
      RECT 1.975000  2.175000 2.165000 2.635000 ;
      RECT 2.335000  0.085000 2.665000 0.595000 ;
      RECT 2.335000  2.005000 2.665000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__a21boi_0
MACRO sky130_fd_sc_hd__a21boi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.760000 0.995000 2.155000 1.345000 ;
        RECT 1.945000 0.375000 2.155000 0.995000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.350000 0.995000 2.640000 1.345000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.975000 0.335000 1.665000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.551000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.045000 1.580000 1.345000 ;
        RECT 1.045000 1.345000 1.375000 2.455000 ;
        RECT 1.335000 0.265000 1.765000 0.795000 ;
        RECT 1.335000 0.795000 1.580000 1.045000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.095000  1.845000 0.855000 2.045000 ;
      RECT 0.095000  2.045000 0.355000 2.435000 ;
      RECT 0.365000  0.265000 0.745000 0.715000 ;
      RECT 0.515000  0.715000 0.745000 1.165000 ;
      RECT 0.515000  1.165000 0.855000 1.845000 ;
      RECT 0.525000  2.225000 0.855000 2.635000 ;
      RECT 0.925000  0.085000 1.155000 0.865000 ;
      RECT 1.545000  1.525000 2.585000 1.725000 ;
      RECT 1.545000  1.725000 1.735000 2.455000 ;
      RECT 1.905000  1.905000 2.235000 2.635000 ;
      RECT 2.325000  0.085000 2.655000 0.815000 ;
      RECT 2.415000  1.725000 2.585000 2.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__a21boi_1
MACRO sky130_fd_sc_hd__einvn_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 0.765000 1.755000 1.955000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.650000 1.725000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.275600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.160000 0.255000 1.755000 0.595000 ;
        RECT 1.160000 0.595000 1.330000 2.125000 ;
        RECT 1.160000 2.125000 1.755000 2.465000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.085000  0.255000 0.360000 0.655000 ;
      RECT 0.085000  0.655000 0.990000 0.825000 ;
      RECT 0.085000  1.895000 0.990000 2.065000 ;
      RECT 0.085000  2.065000 0.400000 2.465000 ;
      RECT 0.530000  0.085000 0.990000 0.485000 ;
      RECT 0.570000  2.235000 0.990000 2.635000 ;
      RECT 0.820000  0.825000 0.990000 1.895000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__einvn_0
MACRO sky130_fd_sc_hd__einvn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 0.765000 2.215000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.309000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.510000 1.725000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 1.785000 2.215000 2.465000 ;
        RECT 1.620000 0.255000 2.215000 0.595000 ;
        RECT 1.620000 0.595000 1.800000 1.785000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.255000 0.370000 0.615000 ;
      RECT 0.085000  0.615000 1.450000 0.785000 ;
      RECT 0.085000  1.895000 0.870000 2.065000 ;
      RECT 0.085000  2.065000 0.370000 2.465000 ;
      RECT 0.540000  0.085000 1.440000 0.445000 ;
      RECT 0.540000  2.235000 0.870000 2.635000 ;
      RECT 0.685000  0.785000 1.450000 1.615000 ;
      RECT 0.685000  1.615000 0.870000 1.895000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__einvn_1
MACRO sky130_fd_sc_hd__einvn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.645000 0.995000 7.800000 1.285000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.375500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.345000 1.325000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.870000 0.620000 8.195000 0.825000 ;
        RECT 4.870000 1.455000 8.195000 1.625000 ;
        RECT 4.870000 1.625000 5.200000 2.125000 ;
        RECT 5.710000 1.625000 6.040000 2.125000 ;
        RECT 6.550000 1.625000 6.880000 2.125000 ;
        RECT 7.390000 1.625000 7.720000 2.125000 ;
        RECT 7.970000 0.825000 8.195000 1.455000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.090000  0.255000 0.345000 0.655000 ;
      RECT 0.090000  0.655000 0.845000 0.825000 ;
      RECT 0.090000  1.495000 0.845000 1.665000 ;
      RECT 0.090000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  0.825000 0.845000 0.995000 ;
      RECT 0.515000  0.995000 4.475000 1.325000 ;
      RECT 0.515000  1.325000 0.845000 1.495000 ;
      RECT 0.515000  1.835000 0.845000 2.635000 ;
      RECT 1.015000  0.255000 1.285000 0.655000 ;
      RECT 1.015000  0.655000 4.700000 0.825000 ;
      RECT 1.015000  1.495000 4.700000 1.665000 ;
      RECT 1.015000  1.665000 1.240000 2.465000 ;
      RECT 1.410000  1.835000 1.740000 2.635000 ;
      RECT 1.455000  0.085000 1.785000 0.485000 ;
      RECT 1.910000  1.665000 2.080000 2.465000 ;
      RECT 1.955000  0.255000 2.125000 0.655000 ;
      RECT 2.250000  1.835000 2.580000 2.635000 ;
      RECT 2.295000  0.085000 2.625000 0.485000 ;
      RECT 2.750000  1.665000 2.920000 2.465000 ;
      RECT 2.795000  0.255000 2.965000 0.655000 ;
      RECT 3.090000  1.835000 3.420000 2.635000 ;
      RECT 3.135000  0.085000 3.465000 0.485000 ;
      RECT 3.590000  1.665000 3.760000 2.465000 ;
      RECT 3.635000  0.255000 3.805000 0.655000 ;
      RECT 3.930000  1.835000 4.280000 2.635000 ;
      RECT 3.975000  0.085000 4.315000 0.485000 ;
      RECT 4.450000  1.665000 4.700000 2.295000 ;
      RECT 4.450000  2.295000 8.195000 2.465000 ;
      RECT 4.485000  0.255000 8.195000 0.450000 ;
      RECT 4.485000  0.450000 4.700000 0.655000 ;
      RECT 5.370000  1.795000 5.540000 2.295000 ;
      RECT 6.210000  1.795000 6.380000 2.295000 ;
      RECT 7.050000  1.795000 7.220000 2.295000 ;
      RECT 7.890000  1.795000 8.195000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
END sky130_fd_sc_hd__einvn_8
MACRO sky130_fd_sc_hd__einvn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 1.075000 3.135000 1.275000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.441000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.325000 1.385000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.694800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.445000 3.135000 1.695000 ;
        RECT 2.365000 0.595000 2.695000 0.845000 ;
        RECT 2.365000 0.845000 2.615000 1.445000 ;
        RECT 2.785000 1.695000 3.135000 2.465000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.840000 0.825000 ;
      RECT 0.085000  1.555000 0.895000 1.725000 ;
      RECT 0.085000  1.725000 0.345000 2.465000 ;
      RECT 0.495000  0.825000 0.840000 0.995000 ;
      RECT 0.495000  0.995000 2.035000 1.275000 ;
      RECT 0.495000  1.275000 0.895000 1.555000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  1.895000 0.895000 2.635000 ;
      RECT 1.015000  0.255000 1.280000 0.655000 ;
      RECT 1.015000  0.655000 2.195000 0.825000 ;
      RECT 1.070000  1.445000 1.775000 1.865000 ;
      RECT 1.070000  1.865000 2.615000 2.085000 ;
      RECT 1.070000  2.085000 1.240000 2.465000 ;
      RECT 1.410000  2.255000 2.275000 2.635000 ;
      RECT 1.450000  0.085000 1.780000 0.485000 ;
      RECT 1.950000  0.255000 3.135000 0.425000 ;
      RECT 1.950000  0.425000 2.195000 0.655000 ;
      RECT 2.445000  2.085000 2.615000 2.465000 ;
      RECT 2.865000  0.425000 3.135000 0.775000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__einvn_2
MACRO sky130_fd_sc_hd__einvn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.530000 0.620000 4.975000 1.325000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.811500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.345000 1.325000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.190000 0.620000 4.360000 1.480000 ;
        RECT 3.190000 1.480000 3.520000 2.075000 ;
        RECT 4.030000 1.480000 4.360000 2.075000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.655000 ;
      RECT 0.085000  0.655000 0.845000 0.825000 ;
      RECT 0.085000  1.495000 0.845000 1.665000 ;
      RECT 0.085000  1.665000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.485000 ;
      RECT 0.515000  0.825000 0.845000 0.995000 ;
      RECT 0.515000  0.995000 3.020000 1.325000 ;
      RECT 0.515000  1.325000 0.845000 1.495000 ;
      RECT 0.515000  1.835000 0.845000 2.635000 ;
      RECT 1.015000  0.255000 1.285000 0.655000 ;
      RECT 1.015000  0.655000 2.995000 0.825000 ;
      RECT 1.015000  1.495000 3.020000 1.665000 ;
      RECT 1.015000  1.665000 1.240000 2.465000 ;
      RECT 1.410000  1.835000 1.740000 2.635000 ;
      RECT 1.455000  0.085000 1.785000 0.485000 ;
      RECT 1.910000  1.665000 2.080000 2.465000 ;
      RECT 1.955000  0.255000 2.125000 0.655000 ;
      RECT 2.250000  1.835000 2.640000 2.635000 ;
      RECT 2.295000  0.085000 2.625000 0.485000 ;
      RECT 2.810000  1.665000 3.020000 2.295000 ;
      RECT 2.810000  2.295000 4.975000 2.465000 ;
      RECT 2.825000  0.255000 4.975000 0.450000 ;
      RECT 2.825000  0.450000 2.995000 0.655000 ;
      RECT 3.690000  1.650000 3.860000 2.295000 ;
      RECT 4.530000  1.650000 4.975000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__einvn_4
MACRO sky130_fd_sc_hd__o221a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.075000 3.605000 1.445000 ;
        RECT 3.005000 1.445000 4.775000 1.615000 ;
        RECT 4.525000 1.075000 5.035000 1.275000 ;
        RECT 4.525000 1.275000 4.775000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775000 1.075000 4.355000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.075000 1.520000 1.445000 ;
        RECT 1.025000 1.445000 2.745000 1.615000 ;
        RECT 2.415000 1.075000 2.745000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.690000 1.075000 2.245000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.440000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235000 0.255000 5.565000 0.725000 ;
        RECT 5.235000 0.725000 6.405000 0.735000 ;
        RECT 5.235000 0.735000 6.920000 0.905000 ;
        RECT 5.315000 1.785000 5.900000 1.955000 ;
        RECT 5.315000 1.955000 5.525000 2.465000 ;
        RECT 5.730000 1.445000 6.920000 1.615000 ;
        RECT 5.730000 1.615000 5.900000 1.785000 ;
        RECT 6.075000 0.255000 6.405000 0.725000 ;
        RECT 6.115000 1.615000 6.365000 2.465000 ;
        RECT 6.575000 0.905000 6.920000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.085000  0.255000 2.955000 0.475000 ;
      RECT 0.085000  0.475000 0.345000 0.895000 ;
      RECT 0.145000  1.455000 0.395000 2.635000 ;
      RECT 0.515000  0.645000 0.845000 0.865000 ;
      RECT 0.565000  1.445000 0.845000 1.785000 ;
      RECT 0.565000  1.785000 5.145000 1.955000 ;
      RECT 0.565000  1.955000 0.815000 2.465000 ;
      RECT 0.610000  0.865000 0.845000 1.445000 ;
      RECT 0.985000  2.125000 1.235000 2.635000 ;
      RECT 1.015000  0.475000 1.185000 0.905000 ;
      RECT 1.355000  0.645000 2.535000 0.715000 ;
      RECT 1.355000  0.715000 3.885000 0.725000 ;
      RECT 1.355000  0.725000 4.725000 0.905000 ;
      RECT 1.405000  2.125000 1.655000 2.295000 ;
      RECT 1.405000  2.295000 2.495000 2.465000 ;
      RECT 1.825000  1.955000 2.075000 2.125000 ;
      RECT 2.245000  2.125000 2.495000 2.295000 ;
      RECT 2.665000  2.125000 3.425000 2.635000 ;
      RECT 3.145000  0.085000 3.385000 0.545000 ;
      RECT 3.555000  0.255000 3.885000 0.715000 ;
      RECT 3.595000  2.125000 3.845000 2.295000 ;
      RECT 3.595000  2.295000 4.685000 2.465000 ;
      RECT 4.015000  1.955000 4.265000 2.125000 ;
      RECT 4.055000  0.085000 4.225000 0.555000 ;
      RECT 4.395000  0.255000 4.725000 0.725000 ;
      RECT 4.435000  2.125000 4.685000 2.295000 ;
      RECT 4.855000  2.125000 5.105000 2.635000 ;
      RECT 4.895000  0.085000 5.065000 0.905000 ;
      RECT 4.975000  1.445000 5.375000 1.615000 ;
      RECT 4.975000  1.615000 5.145000 1.785000 ;
      RECT 5.205000  1.075000 6.405000 1.275000 ;
      RECT 5.205000  1.275000 5.375000 1.445000 ;
      RECT 5.695000  2.125000 5.945000 2.635000 ;
      RECT 5.735000  0.085000 5.905000 0.555000 ;
      RECT 6.535000  1.795000 6.785000 2.635000 ;
      RECT 6.575000  0.085000 6.830000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__o221a_4
MACRO sky130_fd_sc_hd__o221a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.680000 1.075000 3.130000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 1.075000 2.490000 1.285000 ;
        RECT 2.005000 1.285000 2.380000 1.705000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.925000 1.075000 1.255000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 1.075000 1.815000 1.325000 ;
        RECT 1.495000 1.325000 1.815000 1.705000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.415000 1.285000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.370000 0.265000 4.055000 0.905000 ;
        RECT 3.390000 1.875000 4.055000 2.465000 ;
        RECT 3.805000 0.905000 4.055000 1.875000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.240000  1.455000 1.325000 1.625000 ;
      RECT 0.240000  1.625000 0.540000 2.465000 ;
      RECT 0.245000  0.255000 0.575000 0.645000 ;
      RECT 0.245000  0.645000 0.755000 0.825000 ;
      RECT 0.585000  0.825000 0.755000 1.455000 ;
      RECT 0.735000  1.795000 0.985000 2.635000 ;
      RECT 0.745000  0.305000 1.930000 0.475000 ;
      RECT 1.155000  1.625000 1.325000 1.875000 ;
      RECT 1.155000  1.875000 2.720000 2.045000 ;
      RECT 1.160000  0.645000 1.545000 0.735000 ;
      RECT 1.160000  0.735000 2.860000 0.905000 ;
      RECT 1.575000  2.045000 2.380000 2.465000 ;
      RECT 2.190000  0.085000 2.360000 0.555000 ;
      RECT 2.530000  0.270000 2.860000 0.735000 ;
      RECT 2.550000  1.455000 3.470000 1.625000 ;
      RECT 2.550000  1.625000 2.720000 1.875000 ;
      RECT 2.890000  1.795000 3.220000 2.635000 ;
      RECT 3.030000  0.085000 3.200000 0.905000 ;
      RECT 3.300000  1.075000 3.635000 1.285000 ;
      RECT 3.300000  1.285000 3.470000 1.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o221a_1
MACRO sky130_fd_sc_hd__o221a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.635000 1.075000 3.075000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.980000 1.075000 2.465000 1.285000 ;
        RECT 1.980000 1.285000 2.285000 1.705000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885000 1.075000 1.230000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.400000 1.075000 1.790000 1.275000 ;
        RECT 1.500000 1.275000 1.790000 1.705000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.345000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.295000 0.265000 3.625000 0.735000 ;
        RECT 3.295000 0.735000 4.055000 0.905000 ;
        RECT 3.295000 1.875000 4.055000 2.045000 ;
        RECT 3.295000 2.045000 3.545000 2.465000 ;
        RECT 3.745000 0.905000 4.055000 1.875000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120000 -0.085000 0.290000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.170000  0.255000 0.500000 0.635000 ;
      RECT 0.170000  0.635000 0.715000 0.805000 ;
      RECT 0.250000  1.495000 1.330000 1.670000 ;
      RECT 0.250000  1.670000 0.580000 2.465000 ;
      RECT 0.545000  0.805000 0.715000 1.445000 ;
      RECT 0.545000  1.445000 1.330000 1.495000 ;
      RECT 0.670000  0.295000 1.855000 0.465000 ;
      RECT 0.750000  1.850000 0.990000 2.635000 ;
      RECT 1.085000  0.645000 1.470000 0.735000 ;
      RECT 1.085000  0.735000 2.785000 0.905000 ;
      RECT 1.160000  1.670000 1.330000 1.875000 ;
      RECT 1.160000  1.875000 2.625000 2.045000 ;
      RECT 1.550000  2.045000 2.305000 2.465000 ;
      RECT 2.115000  0.085000 2.285000 0.555000 ;
      RECT 2.455000  0.270000 2.785000 0.735000 ;
      RECT 2.455000  1.455000 3.415000 1.625000 ;
      RECT 2.455000  1.625000 2.625000 1.875000 ;
      RECT 2.795000  1.795000 3.125000 2.635000 ;
      RECT 2.955000  0.085000 3.125000 0.905000 ;
      RECT 3.245000  1.075000 3.575000 1.285000 ;
      RECT 3.245000  1.285000 3.415000 1.455000 ;
      RECT 3.715000  2.215000 4.055000 2.635000 ;
      RECT 3.795000  0.085000 3.965000 0.565000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__o221a_2
MACRO sky130_fd_sc_hd__dfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.160000 0.265000 9.495000 1.695000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.030000 1.535000 10.420000 2.080000 ;
        RECT 10.040000 0.310000 10.420000 0.825000 ;
        RECT 10.120000 2.080000 10.420000 2.465000 ;
        RECT 10.250000 0.825000 10.420000 1.535000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.090000  0.345000  0.345000 0.635000 ;
      RECT  0.090000  0.635000  0.840000 0.805000 ;
      RECT  0.090000  1.795000  0.840000 1.965000 ;
      RECT  0.090000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.610000  0.805000  0.840000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.545000  0.085000  1.875000 0.445000 ;
      RECT  1.850000  2.175000  2.100000 2.635000 ;
      RECT  2.045000  0.305000  2.540000 0.475000 ;
      RECT  2.045000  0.475000  2.215000 1.835000 ;
      RECT  2.045000  1.835000  2.440000 2.005000 ;
      RECT  2.270000  2.005000  2.440000 2.135000 ;
      RECT  2.270000  2.135000  2.520000 2.465000 ;
      RECT  2.385000  0.765000  2.735000 1.385000 ;
      RECT  2.610000  1.575000  3.075000 1.965000 ;
      RECT  2.735000  2.135000  3.415000 2.465000 ;
      RECT  2.745000  0.305000  3.600000 0.475000 ;
      RECT  2.905000  0.765000  3.260000 0.985000 ;
      RECT  2.905000  0.985000  3.075000 1.575000 ;
      RECT  3.245000  1.185000  4.935000 1.355000 ;
      RECT  3.245000  1.355000  3.415000 2.135000 ;
      RECT  3.430000  0.475000  3.600000 1.185000 ;
      RECT  3.585000  1.865000  4.660000 2.035000 ;
      RECT  3.585000  2.035000  3.755000 2.375000 ;
      RECT  3.775000  1.525000  5.275000 1.695000 ;
      RECT  3.990000  2.205000  4.320000 2.635000 ;
      RECT  4.475000  0.085000  4.805000 0.545000 ;
      RECT  4.490000  2.035000  4.660000 2.375000 ;
      RECT  4.765000  1.005000  4.935000 1.185000 ;
      RECT  4.955000  2.175000  5.325000 2.635000 ;
      RECT  5.015000  0.275000  5.365000 0.445000 ;
      RECT  5.015000  0.445000  5.275000 0.835000 ;
      RECT  5.105000  0.835000  5.275000 1.525000 ;
      RECT  5.105000  1.695000  5.275000 1.835000 ;
      RECT  5.105000  1.835000  5.665000 2.005000 ;
      RECT  5.465000  0.705000  5.675000 1.495000 ;
      RECT  5.465000  1.495000  6.140000 1.655000 ;
      RECT  5.465000  1.655000  6.430000 1.665000 ;
      RECT  5.495000  2.005000  5.665000 2.465000 ;
      RECT  5.585000  0.255000  6.535000 0.535000 ;
      RECT  5.845000  0.705000  6.195000 1.325000 ;
      RECT  5.900000  2.125000  6.770000 2.465000 ;
      RECT  5.970000  1.665000  6.430000 1.955000 ;
      RECT  6.365000  0.535000  6.535000 1.315000 ;
      RECT  6.365000  1.315000  6.770000 1.485000 ;
      RECT  6.600000  1.485000  6.770000 1.575000 ;
      RECT  6.600000  1.575000  7.820000 1.745000 ;
      RECT  6.600000  1.745000  6.770000 2.125000 ;
      RECT  6.705000  0.085000  6.895000 0.525000 ;
      RECT  6.705000  0.695000  7.235000 0.865000 ;
      RECT  6.705000  0.865000  6.925000 1.145000 ;
      RECT  6.940000  2.175000  7.190000 2.635000 ;
      RECT  7.065000  0.295000  7.985000 0.465000 ;
      RECT  7.065000  0.465000  7.235000 0.695000 ;
      RECT  7.360000  1.915000  8.160000 2.085000 ;
      RECT  7.360000  2.085000  7.530000 2.375000 ;
      RECT  7.710000  2.255000  8.055000 2.635000 ;
      RECT  7.815000  0.465000  7.985000 0.995000 ;
      RECT  7.815000  0.995000  8.160000 1.075000 ;
      RECT  7.815000  1.075000  8.650000 1.295000 ;
      RECT  7.990000  1.295000  8.650000 1.325000 ;
      RECT  7.990000  1.325000  8.160000 1.915000 ;
      RECT  8.335000  0.345000  8.585000 0.715000 ;
      RECT  8.335000  0.715000  8.990000 0.885000 ;
      RECT  8.335000  1.795000  8.990000 1.865000 ;
      RECT  8.335000  1.865000  9.835000 2.035000 ;
      RECT  8.335000  2.035000  8.560000 2.465000 ;
      RECT  8.730000  2.205000  9.070000 2.635000 ;
      RECT  8.755000  0.085000  8.990000 0.545000 ;
      RECT  8.820000  0.885000  8.990000 1.795000 ;
      RECT  9.620000  2.255000  9.950000 2.635000 ;
      RECT  9.665000  0.995000 10.080000 1.325000 ;
      RECT  9.665000  1.325000  9.835000 1.865000 ;
      RECT  9.700000  0.085000  9.870000 0.825000 ;
      RECT 10.590000  0.085000 10.760000 0.930000 ;
      RECT 10.590000  1.445000 10.760000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.610000  1.105000  0.780000 1.275000 ;
      RECT  1.015000  1.785000  1.185000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.105000  2.615000 1.275000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  1.785000  3.075000 1.955000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.025000  1.105000  6.195000 1.275000 ;
      RECT  6.025000  1.785000  6.195000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.075000 0.840000 1.120000 ;
      RECT 0.550000 1.120000 6.255000 1.260000 ;
      RECT 0.550000 1.260000 0.840000 1.305000 ;
      RECT 0.955000 1.755000 1.245000 1.800000 ;
      RECT 0.955000 1.800000 6.255000 1.940000 ;
      RECT 0.955000 1.940000 1.245000 1.985000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrbp_2
MACRO sky130_fd_sc_hd__dfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.600000 1.455000 9.005000 2.465000 ;
        RECT 8.675000 0.275000 9.005000 1.455000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.180000 0.265000 10.435000 0.795000 ;
        RECT 10.180000 1.445000 10.435000 2.325000 ;
        RECT 10.225000 0.795000 10.435000 1.445000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.770000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.580000 0.085000 ;
      RECT 0.000000  2.635000 10.580000 2.805000 ;
      RECT 0.090000  0.345000  0.345000 0.635000 ;
      RECT 0.090000  0.635000  0.840000 0.805000 ;
      RECT 0.090000  1.795000  0.840000 1.965000 ;
      RECT 0.090000  1.965000  0.345000 2.465000 ;
      RECT 0.515000  0.085000  0.845000 0.465000 ;
      RECT 0.515000  2.135000  0.845000 2.635000 ;
      RECT 0.610000  0.805000  0.840000 1.795000 ;
      RECT 1.015000  0.345000  1.185000 2.465000 ;
      RECT 1.545000  0.085000  1.875000 0.445000 ;
      RECT 1.850000  2.175000  2.100000 2.635000 ;
      RECT 2.045000  0.305000  2.540000 0.475000 ;
      RECT 2.045000  0.475000  2.215000 1.835000 ;
      RECT 2.045000  1.835000  2.440000 2.005000 ;
      RECT 2.270000  2.005000  2.440000 2.135000 ;
      RECT 2.270000  2.135000  2.520000 2.465000 ;
      RECT 2.385000  0.765000  2.735000 1.385000 ;
      RECT 2.610000  1.575000  3.075000 1.965000 ;
      RECT 2.735000  2.135000  3.415000 2.465000 ;
      RECT 2.745000  0.305000  3.600000 0.475000 ;
      RECT 2.905000  0.765000  3.260000 0.985000 ;
      RECT 2.905000  0.985000  3.075000 1.575000 ;
      RECT 3.245000  1.185000  4.935000 1.355000 ;
      RECT 3.245000  1.355000  3.415000 2.135000 ;
      RECT 3.430000  0.475000  3.600000 1.185000 ;
      RECT 3.585000  1.865000  4.660000 2.035000 ;
      RECT 3.585000  2.035000  3.755000 2.375000 ;
      RECT 3.775000  1.525000  5.275000 1.695000 ;
      RECT 3.990000  2.205000  4.320000 2.635000 ;
      RECT 4.475000  0.085000  4.805000 0.545000 ;
      RECT 4.490000  2.035000  4.660000 2.375000 ;
      RECT 4.765000  1.005000  4.935000 1.185000 ;
      RECT 4.955000  2.175000  5.325000 2.635000 ;
      RECT 5.015000  0.275000  5.365000 0.445000 ;
      RECT 5.015000  0.445000  5.275000 0.835000 ;
      RECT 5.105000  0.835000  5.275000 1.525000 ;
      RECT 5.105000  1.695000  5.275000 1.835000 ;
      RECT 5.105000  1.835000  5.665000 2.005000 ;
      RECT 5.465000  0.705000  5.675000 1.495000 ;
      RECT 5.465000  1.495000  6.140000 1.655000 ;
      RECT 5.465000  1.655000  6.430000 1.665000 ;
      RECT 5.495000  2.005000  5.665000 2.465000 ;
      RECT 5.585000  0.255000  6.535000 0.535000 ;
      RECT 5.845000  0.705000  6.195000 1.325000 ;
      RECT 5.900000  2.125000  6.770000 2.465000 ;
      RECT 5.970000  1.665000  6.430000 1.955000 ;
      RECT 6.365000  0.535000  6.535000 1.315000 ;
      RECT 6.365000  1.315000  6.770000 1.485000 ;
      RECT 6.600000  1.485000  6.770000 1.575000 ;
      RECT 6.600000  1.575000  7.820000 1.745000 ;
      RECT 6.600000  1.745000  6.770000 2.125000 ;
      RECT 6.705000  0.085000  6.895000 0.525000 ;
      RECT 6.705000  0.695000  7.235000 0.865000 ;
      RECT 6.705000  0.865000  6.925000 1.145000 ;
      RECT 6.940000  2.175000  7.190000 2.635000 ;
      RECT 7.065000  0.295000  8.135000 0.465000 ;
      RECT 7.065000  0.465000  7.235000 0.695000 ;
      RECT 7.360000  1.915000  8.160000 2.085000 ;
      RECT 7.360000  2.085000  7.530000 2.375000 ;
      RECT 7.710000  2.255000  8.430000 2.635000 ;
      RECT 7.815000  0.465000  8.135000 0.820000 ;
      RECT 7.815000  0.820000  8.140000 0.995000 ;
      RECT 7.815000  0.995000  8.435000 1.295000 ;
      RECT 7.990000  1.295000  8.435000 1.325000 ;
      RECT 7.990000  1.325000  8.160000 1.915000 ;
      RECT 8.335000  0.085000  8.505000 0.770000 ;
      RECT 9.195000  0.345000  9.445000 0.995000 ;
      RECT 9.195000  0.995000 10.055000 1.325000 ;
      RECT 9.195000  1.325000  9.525000 2.425000 ;
      RECT 9.760000  0.085000  9.930000 0.680000 ;
      RECT 9.760000  1.495000  9.930000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.610000  1.105000  0.780000 1.275000 ;
      RECT  1.015000  1.785000  1.185000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  1.105000  2.615000 1.275000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  1.785000  3.075000 1.955000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.025000  1.105000  6.195000 1.275000 ;
      RECT  6.025000  1.785000  6.195000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.075000 0.840000 1.120000 ;
      RECT 0.550000 1.120000 6.255000 1.260000 ;
      RECT 0.550000 1.260000 0.840000 1.305000 ;
      RECT 0.955000 1.755000 1.245000 1.800000 ;
      RECT 0.955000 1.800000 6.255000 1.940000 ;
      RECT 0.955000 1.940000 1.245000 1.985000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrbp_1
MACRO sky130_fd_sc_hd__a211o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.035000 1.020000 5.380000 1.330000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.495000 1.020000 4.825000 1.510000 ;
        RECT 4.495000 1.510000 5.845000 1.700000 ;
        RECT 5.635000 1.020000 6.225000 1.320000 ;
        RECT 5.635000 1.320000 5.845000 1.510000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.540000 0.985000 2.805000 1.325000 ;
        RECT 2.625000 1.325000 2.805000 1.445000 ;
        RECT 2.625000 1.445000 4.175000 1.700000 ;
        RECT 3.845000 0.985000 4.175000 1.445000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.975000 0.985000 3.645000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.933750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.635000 2.025000 0.875000 ;
        RECT 0.085000 0.875000 0.340000 1.495000 ;
        RECT 0.085000 1.495000 1.640000 1.705000 ;
        RECT 0.595000 1.705000 0.780000 2.465000 ;
        RECT 0.985000 0.255000 1.175000 0.615000 ;
        RECT 0.985000 0.615000 2.025000 0.635000 ;
        RECT 1.450000 1.705000 1.640000 2.465000 ;
        RECT 1.845000 0.255000 2.025000 0.615000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.090000  1.875000 0.425000 2.635000 ;
      RECT 0.485000  0.085000 0.815000 0.465000 ;
      RECT 0.525000  1.045000 2.370000 1.325000 ;
      RECT 0.950000  1.875000 1.280000 2.635000 ;
      RECT 1.345000  0.085000 1.675000 0.445000 ;
      RECT 1.810000  1.835000 2.060000 2.635000 ;
      RECT 2.185000  1.325000 2.370000 1.505000 ;
      RECT 2.185000  1.505000 2.455000 1.675000 ;
      RECT 2.195000  0.615000 5.490000 0.805000 ;
      RECT 2.195000  0.805000 2.370000 1.045000 ;
      RECT 2.220000  0.085000 2.555000 0.445000 ;
      RECT 2.280000  1.675000 2.455000 1.870000 ;
      RECT 2.280000  1.870000 3.510000 2.040000 ;
      RECT 2.320000  2.210000 4.450000 2.465000 ;
      RECT 2.725000  0.255000 2.970000 0.615000 ;
      RECT 3.140000  0.085000 3.470000 0.445000 ;
      RECT 3.640000  0.255000 4.020000 0.615000 ;
      RECT 4.120000  1.880000 6.345000 2.105000 ;
      RECT 4.120000  2.105000 4.450000 2.210000 ;
      RECT 4.190000  0.085000 4.560000 0.445000 ;
      RECT 4.620000  2.275000 4.950000 2.635000 ;
      RECT 5.160000  0.275000 5.490000 0.615000 ;
      RECT 5.160000  2.105000 5.420000 2.465000 ;
      RECT 5.590000  2.275000 5.920000 2.635000 ;
      RECT 6.015000  0.085000 6.345000 0.805000 ;
      RECT 6.015000  1.535000 6.345000 1.880000 ;
      RECT 6.090000  2.105000 6.345000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
END sky130_fd_sc_hd__a211o_4
MACRO sky130_fd_sc_hd__a211o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 0.995000 2.060000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 0.995000 1.305000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.240000 0.995000 2.675000 1.325000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855000 0.995000 3.125000 1.325000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.437250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.265000 0.425000 1.685000 ;
        RECT 0.090000 1.685000 0.355000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.135000 -0.085000 0.305000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.525000  1.915000 0.855000 2.635000 ;
      RECT 0.600000  0.625000 3.085000 0.815000 ;
      RECT 0.600000  0.815000 0.825000 1.505000 ;
      RECT 0.600000  1.505000 3.095000 1.685000 ;
      RECT 0.605000  0.085000 1.350000 0.455000 ;
      RECT 1.045000  1.865000 2.235000 2.095000 ;
      RECT 1.045000  2.095000 1.305000 2.455000 ;
      RECT 1.475000  2.265000 1.805000 2.635000 ;
      RECT 1.915000  0.265000 2.170000 0.625000 ;
      RECT 1.975000  2.095000 2.235000 2.455000 ;
      RECT 2.350000  0.085000 2.680000 0.455000 ;
      RECT 2.805000  1.685000 3.095000 2.455000 ;
      RECT 2.860000  0.265000 3.085000 0.625000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a211o_1
MACRO sky130_fd_sc_hd__a211o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.980000 1.045000 2.450000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.480000 1.045000 1.810000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.620000 1.045000 3.070000 1.275000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.260000 1.045000 3.595000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.452000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.255000 0.775000 0.635000 ;
        RECT 0.555000 0.635000 0.785000 2.335000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.085000 0.385000 0.905000 ;
      RECT 0.090000  1.490000 0.385000 2.635000 ;
      RECT 0.945000  0.085000 1.795000 0.445000 ;
      RECT 1.000000  0.695000 3.585000 0.875000 ;
      RECT 1.000000  0.875000 1.310000 1.490000 ;
      RECT 1.000000  1.490000 3.585000 1.660000 ;
      RECT 1.000000  1.830000 1.255000 2.635000 ;
      RECT 1.455000  1.840000 2.795000 2.020000 ;
      RECT 1.455000  2.020000 1.785000 2.465000 ;
      RECT 1.955000  2.190000 2.230000 2.635000 ;
      RECT 2.275000  0.275000 2.605000 0.695000 ;
      RECT 2.465000  2.020000 2.795000 2.465000 ;
      RECT 2.810000  0.085000 3.085000 0.525000 ;
      RECT 3.255000  0.275000 3.585000 0.695000 ;
      RECT 3.255000  1.660000 3.585000 2.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a211o_2
MACRO sky130_fd_sc_hd__and3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.955000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.790000 2.125000 2.265000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.305000 2.185000 0.725000 ;
        RECT 1.985000 0.725000 2.395000 1.245000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.860000 1.765000 3.135000 2.465000 ;
        RECT 2.875000 0.255000 3.135000 0.735000 ;
        RECT 2.965000 0.735000 3.135000 1.765000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.905000 ;
      RECT 0.085000  2.125000 0.345000 2.635000 ;
      RECT 0.515000  0.485000 0.845000 0.905000 ;
      RECT 0.595000  0.905000 0.845000 0.995000 ;
      RECT 0.595000  0.995000 1.390000 1.245000 ;
      RECT 0.595000  1.245000 0.765000 2.465000 ;
      RECT 1.005000  1.425000 2.795000 1.595000 ;
      RECT 1.005000  1.595000 1.255000 1.960000 ;
      RECT 1.005000  2.130000 1.620000 2.635000 ;
      RECT 1.025000  0.305000 1.815000 0.570000 ;
      RECT 1.425000  1.765000 1.755000 1.955000 ;
      RECT 1.425000  1.955000 1.620000 2.130000 ;
      RECT 1.560000  0.570000 1.815000 1.425000 ;
      RECT 1.975000  1.595000 2.690000 1.890000 ;
      RECT 2.375000  0.085000 2.705000 0.545000 ;
      RECT 2.435000  2.090000 2.650000 2.635000 ;
      RECT 2.565000  0.995000 2.795000 1.425000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__and3b_1
MACRO sky130_fd_sc_hd__and3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.715000 0.615000 3.995000 1.705000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 0.725000 1.235000 1.340000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 1.715000 1.340000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.934000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225000 1.535000 3.535000 1.705000 ;
        RECT 2.285000 0.515000 2.475000 0.615000 ;
        RECT 2.285000 0.615000 3.535000 0.845000 ;
        RECT 3.145000 0.255000 3.335000 0.615000 ;
        RECT 3.270000 0.845000 3.535000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.150000  0.255000 0.635000 0.355000 ;
      RECT 0.150000  0.355000 1.600000 0.545000 ;
      RECT 0.150000  0.545000 0.635000 0.805000 ;
      RECT 0.150000  0.805000 0.370000 1.495000 ;
      RECT 0.150000  1.495000 0.510000 2.165000 ;
      RECT 0.540000  0.995000 0.850000 1.325000 ;
      RECT 0.680000  1.325000 0.850000 1.875000 ;
      RECT 0.680000  1.875000 4.445000 2.105000 ;
      RECT 0.730000  2.275000 1.180000 2.635000 ;
      RECT 1.280000  1.525000 2.055000 1.695000 ;
      RECT 1.420000  0.545000 1.600000 0.615000 ;
      RECT 1.420000  0.615000 2.115000 0.805000 ;
      RECT 1.745000  2.275000 2.075000 2.635000 ;
      RECT 1.780000  0.085000 2.110000 0.445000 ;
      RECT 1.885000  0.805000 2.115000 1.020000 ;
      RECT 1.885000  1.020000 3.100000 1.355000 ;
      RECT 1.885000  1.355000 2.055000 1.525000 ;
      RECT 2.645000  0.085000 2.975000 0.445000 ;
      RECT 2.645000  2.275000 2.980000 2.635000 ;
      RECT 3.505000  0.085000 3.835000 0.445000 ;
      RECT 3.505000  2.275000 3.835000 2.635000 ;
      RECT 4.165000  0.425000 4.445000 1.875000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__and3b_4
MACRO sky130_fd_sc_hd__and3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.745000 0.410000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.815000 2.125000 2.290000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.010000 0.305000 2.220000 0.765000 ;
        RECT 2.010000 0.765000 2.420000 1.245000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875000 1.795000 3.160000 2.465000 ;
        RECT 2.915000 0.255000 3.160000 0.715000 ;
        RECT 2.990000 0.715000 3.160000 0.925000 ;
        RECT 2.990000 0.925000 3.595000 1.445000 ;
        RECT 2.990000 1.445000 3.160000 1.795000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 0.355000 0.575000 ;
      RECT 0.085000  1.575000 0.400000 2.635000 ;
      RECT 0.580000  0.305000 0.855000 1.015000 ;
      RECT 0.580000  1.015000 1.415000 1.245000 ;
      RECT 0.580000  1.245000 0.855000 1.905000 ;
      RECT 1.030000  2.130000 1.645000 2.635000 ;
      RECT 1.050000  1.425000 2.820000 1.595000 ;
      RECT 1.050000  1.595000 1.285000 1.960000 ;
      RECT 1.055000  0.305000 1.840000 0.570000 ;
      RECT 1.455000  1.765000 1.785000 1.955000 ;
      RECT 1.455000  1.955000 1.645000 2.130000 ;
      RECT 1.585000  0.570000 1.840000 1.425000 ;
      RECT 2.010000  1.595000 2.200000 1.890000 ;
      RECT 2.410000  0.085000 2.740000 0.580000 ;
      RECT 2.460000  1.790000 2.675000 2.635000 ;
      RECT 2.590000  0.995000 2.820000 1.425000 ;
      RECT 3.330000  0.085000 3.595000 0.745000 ;
      RECT 3.330000  1.625000 3.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__and3b_2
MACRO sky130_fd_sc_hd__o21ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.995000 0.410000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.590000 0.995000 0.975000 1.325000 ;
        RECT 0.590000 1.325000 0.785000 2.375000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.202500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.295000 1.750000 1.655000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.517000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.505000 1.315000 1.785000 ;
        RECT 0.965000 1.785000 1.295000 2.465000 ;
        RECT 1.145000 0.955000 1.665000 1.125000 ;
        RECT 1.145000 1.125000 1.315000 1.505000 ;
        RECT 1.495000 0.390000 1.665000 0.955000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.090000  0.265000 0.380000 0.615000 ;
      RECT 0.090000  0.615000 1.305000 0.785000 ;
      RECT 0.090000  1.495000 0.410000 2.635000 ;
      RECT 0.575000  0.085000 0.905000 0.445000 ;
      RECT 1.075000  0.310000 1.305000 0.615000 ;
      RECT 1.495000  1.835000 1.750000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ai_1
MACRO sky130_fd_sc_hd__o21ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 1.055000 0.450000 1.445000 ;
        RECT 0.120000 1.445000 2.095000 1.615000 ;
        RECT 1.600000 1.075000 2.095000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.620000 1.075000 1.420000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815000 0.765000 3.130000 1.400000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.742000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.785000 2.645000 1.965000 ;
        RECT 0.995000 1.965000 1.295000 2.125000 ;
        RECT 2.410000 1.965000 2.645000 2.465000 ;
        RECT 2.435000 0.595000 2.645000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140000 -0.085000 0.310000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.105000  0.255000 0.435000 0.715000 ;
      RECT 0.105000  0.715000 2.265000 0.885000 ;
      RECT 0.105000  1.785000 0.435000 2.635000 ;
      RECT 0.605000  1.785000 0.825000 2.295000 ;
      RECT 0.605000  2.295000 1.715000 2.465000 ;
      RECT 0.615000  0.085000 0.785000 0.545000 ;
      RECT 0.965000  0.255000 1.295000 0.715000 ;
      RECT 1.525000  0.085000 1.695000 0.545000 ;
      RECT 1.525000  2.135000 1.715000 2.295000 ;
      RECT 1.910000  2.175000 2.240000 2.635000 ;
      RECT 1.935000  0.255000 3.125000 0.425000 ;
      RECT 1.935000  0.425000 2.265000 0.715000 ;
      RECT 2.815000  0.425000 3.125000 0.595000 ;
      RECT 2.815000  1.570000 3.125000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ai_2
MACRO sky130_fd_sc_hd__o21ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.015000 1.475000 1.320000 ;
        RECT 0.575000 1.320000 1.475000 1.515000 ;
        RECT 0.575000 1.515000 3.695000 1.685000 ;
        RECT 3.445000 0.990000 3.695000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.070000 3.275000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.905000 1.015000 5.255000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.840000 1.855000 5.150000 2.025000 ;
        RECT 3.935000 1.445000 5.835000 1.700000 ;
        RECT 3.935000 1.700000 5.150000 1.855000 ;
        RECT 4.030000 0.615000 5.835000 0.845000 ;
        RECT 4.080000 2.025000 5.150000 2.085000 ;
        RECT 4.080000 2.085000 4.290000 2.465000 ;
        RECT 4.960000 2.085000 5.150000 2.465000 ;
        RECT 5.425000 0.845000 5.835000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.120000  0.615000 3.860000 0.820000 ;
      RECT 0.120000  1.820000 0.405000 2.635000 ;
      RECT 0.550000  0.085000 0.880000 0.445000 ;
      RECT 0.575000  1.915000 1.670000 2.085000 ;
      RECT 0.575000  2.085000 0.810000 2.465000 ;
      RECT 0.980000  2.255000 1.310000 2.635000 ;
      RECT 1.410000  0.085000 1.740000 0.445000 ;
      RECT 1.480000  2.085000 1.670000 2.275000 ;
      RECT 1.480000  2.275000 3.460000 2.465000 ;
      RECT 2.270000  0.085000 2.600000 0.445000 ;
      RECT 3.130000  0.085000 3.460000 0.445000 ;
      RECT 3.630000  0.255000 5.650000 0.445000 ;
      RECT 3.630000  0.445000 3.860000 0.615000 ;
      RECT 3.630000  2.195000 3.910000 2.635000 ;
      RECT 4.460000  2.255000 4.790000 2.635000 ;
      RECT 5.320000  1.880000 5.650000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ai_4
MACRO sky130_fd_sc_hd__o21ai_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.415000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.100000 1.005000 1.340000 ;
        RECT 0.605000 1.340000 0.775000 1.645000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 1.355000 1.730000 1.685000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.290500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.510000 1.345000 1.680000 ;
        RECT 0.965000 1.680000 1.300000 2.465000 ;
        RECT 1.175000 0.955000 1.740000 1.125000 ;
        RECT 1.175000 1.125000 1.345000 1.510000 ;
        RECT 1.455000 0.280000 1.740000 0.955000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.030000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.120000  0.280000 0.380000 0.615000 ;
      RECT 0.120000  0.615000 1.285000 0.785000 ;
      RECT 0.145000  1.825000 0.475000 2.635000 ;
      RECT 0.550000  0.085000 0.880000 0.445000 ;
      RECT 1.050000  0.280000 1.285000 0.615000 ;
      RECT 1.470000  1.855000 1.725000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__o21ai_0
MACRO sky130_fd_sc_hd__a2111o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.995000 3.290000 1.325000 ;
        RECT 2.985000 0.285000 3.540000 0.845000 ;
        RECT 2.985000 0.845000 3.290000 0.995000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.510000 1.025000 4.010000 1.290000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.400000 0.995000 2.680000 2.465000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.890000 1.050000 2.220000 2.465000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.290000 1.050000 1.720000 1.290000 ;
        RECT 1.515000 1.290000 1.720000 2.465000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.504500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.255000 0.465000 1.620000 ;
        RECT 0.135000 1.620000 0.390000 2.460000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
    PORT
      LAYER pwell ;
        RECT 1.975000 -0.065000 2.145000 0.105000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.565000  1.815000 0.895000 2.635000 ;
      RECT 0.635000  0.085000 1.310000 0.470000 ;
      RECT 0.695000  0.650000 1.915000 0.655000 ;
      RECT 0.695000  0.655000 2.805000 0.825000 ;
      RECT 0.695000  0.825000 0.915000 1.465000 ;
      RECT 0.695000  1.465000 1.345000 1.645000 ;
      RECT 1.135000  1.645000 1.345000 2.460000 ;
      RECT 1.585000  0.260000 1.915000 0.650000 ;
      RECT 2.085000  0.085000 2.430000 0.485000 ;
      RECT 2.600000  0.260000 2.805000 0.655000 ;
      RECT 2.860000  1.495000 3.990000 1.665000 ;
      RECT 2.860000  1.665000 3.145000 2.460000 ;
      RECT 3.325000  1.835000 3.540000 2.635000 ;
      RECT 3.715000  0.085000 3.955000 0.760000 ;
      RECT 3.720000  1.665000 3.990000 2.460000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111o_1
MACRO sky130_fd_sc_hd__a2111o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 0.955000 3.775000 1.740000 ;
        RECT 3.505000 0.290000 3.995000 0.825000 ;
        RECT 3.505000 0.825000 3.775000 0.955000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.945000 0.995000 4.515000 1.740000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.995000 3.195000 1.740000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425000 0.995000 2.735000 2.355000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 0.995000 2.255000 1.325000 ;
        RECT 1.960000 1.325000 2.255000 2.355000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.255000 0.895000 2.390000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.085000 0.435000 0.885000 ;
      RECT 0.085000  1.635000 0.435000 2.635000 ;
      RECT 1.065000  0.085000 2.010000 0.445000 ;
      RECT 1.065000  0.445000 1.325000 0.865000 ;
      RECT 1.065000  1.075000 1.705000 1.325000 ;
      RECT 1.065000  1.495000 1.315000 2.635000 ;
      RECT 1.495000  0.615000 3.335000 0.785000 ;
      RECT 1.495000  0.785000 1.705000 1.075000 ;
      RECT 1.495000  1.325000 1.705000 1.495000 ;
      RECT 1.495000  1.495000 1.785000 2.465000 ;
      RECT 2.180000  0.255000 2.420000 0.615000 ;
      RECT 2.590000  0.085000 2.920000 0.445000 ;
      RECT 3.070000  1.915000 4.515000 2.085000 ;
      RECT 3.070000  2.085000 3.400000 2.465000 ;
      RECT 3.090000  0.255000 3.335000 0.615000 ;
      RECT 3.590000  2.255000 3.920000 2.635000 ;
      RECT 4.090000  2.085000 4.515000 2.465000 ;
      RECT 4.165000  0.085000 4.515000 0.805000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111o_2
MACRO sky130_fd_sc_hd__a2111o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825000 1.075000 4.495000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675000 1.075000 5.625000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.450000 0.975000 3.255000 1.285000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 0.975000 2.280000 1.285000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.370000 1.625000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.165000 0.255000 6.355000 0.635000 ;
        RECT 6.165000 0.635000 7.735000 0.805000 ;
        RECT 6.165000 1.465000 7.735000 1.635000 ;
        RECT 6.165000 1.635000 7.215000 1.715000 ;
        RECT 6.165000 1.715000 6.355000 2.465000 ;
        RECT 7.025000 0.255000 7.215000 0.635000 ;
        RECT 7.025000 1.715000 7.215000 2.465000 ;
        RECT 7.490000 0.805000 7.735000 1.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.110000  1.795000 0.370000 2.295000 ;
      RECT 0.110000  2.295000 2.160000 2.465000 ;
      RECT 0.180000  0.255000 0.440000 0.635000 ;
      RECT 0.180000  0.635000 3.655000 0.805000 ;
      RECT 0.540000  0.805000 0.870000 2.125000 ;
      RECT 0.610000  0.085000 0.940000 0.465000 ;
      RECT 1.040000  1.455000 1.230000 2.295000 ;
      RECT 1.110000  0.255000 1.340000 0.615000 ;
      RECT 1.110000  0.615000 3.655000 0.635000 ;
      RECT 1.400000  1.455000 3.100000 1.625000 ;
      RECT 1.400000  1.625000 1.730000 2.125000 ;
      RECT 1.510000  0.085000 1.840000 0.445000 ;
      RECT 1.900000  1.795000 2.160000 2.295000 ;
      RECT 2.015000  0.255000 2.240000 0.615000 ;
      RECT 2.340000  1.795000 2.675000 2.295000 ;
      RECT 2.340000  2.295000 3.650000 2.465000 ;
      RECT 2.420000  0.085000 3.295000 0.445000 ;
      RECT 2.845000  1.625000 3.100000 2.125000 ;
      RECT 3.320000  1.795000 5.495000 1.995000 ;
      RECT 3.320000  1.995000 3.650000 2.295000 ;
      RECT 3.465000  0.255000 4.585000 0.445000 ;
      RECT 3.465000  0.445000 3.655000 0.615000 ;
      RECT 3.465000  0.805000 3.655000 1.445000 ;
      RECT 3.465000  1.445000 5.975000 1.625000 ;
      RECT 3.825000  0.615000 5.495000 0.785000 ;
      RECT 3.865000  2.165000 4.195000 2.635000 ;
      RECT 4.365000  1.995000 4.625000 2.415000 ;
      RECT 4.805000  0.085000 5.140000 0.445000 ;
      RECT 4.805000  2.255000 5.140000 2.635000 ;
      RECT 5.310000  0.255000 5.495000 0.615000 ;
      RECT 5.310000  1.995000 5.495000 2.465000 ;
      RECT 5.665000  0.085000 5.995000 0.515000 ;
      RECT 5.665000  1.800000 5.995000 2.635000 ;
      RECT 5.795000  1.075000 7.320000 1.245000 ;
      RECT 5.795000  1.245000 5.975000 1.445000 ;
      RECT 6.525000  0.085000 6.855000 0.445000 ;
      RECT 6.525000  1.885000 6.855000 2.635000 ;
      RECT 7.385000  0.085000 7.715000 0.465000 ;
      RECT 7.385000  1.805000 7.715000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__a2111o_4
MACRO sky130_fd_sc_hd__conb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__conb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.605000 1.740000 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.775000 0.915000 1.295000 2.465000 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.275000  1.910000 0.605000 2.635000 ;
      RECT 0.775000  0.085000 1.115000 0.745000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__conb_1
MACRO sky130_fd_sc_hd__or4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.755000 0.995000 2.925000 1.445000 ;
        RECT 2.755000 1.445000 3.190000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195000 0.995000 2.525000 1.450000 ;
        RECT 2.335000 1.450000 2.525000 1.785000 ;
        RECT 2.335000 1.785000 2.635000 2.375000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795000 0.995000 1.965000 1.620000 ;
        RECT 1.795000 1.620000 2.155000 2.375000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.995000 0.445000 1.955000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 1.455000 4.965000 1.625000 ;
        RECT 3.395000 1.625000 3.645000 2.465000 ;
        RECT 3.435000 0.255000 3.685000 0.725000 ;
        RECT 3.435000 0.725000 4.965000 0.905000 ;
        RECT 4.195000 0.255000 4.525000 0.725000 ;
        RECT 4.235000 1.625000 4.485000 2.465000 ;
        RECT 4.725000 0.905000 4.965000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.825000 ;
      RECT 0.085000  2.135000 0.365000 2.635000 ;
      RECT 0.595000  0.435000 0.785000 0.905000 ;
      RECT 0.595000  2.065000 0.785000 2.455000 ;
      RECT 0.615000  0.905000 0.785000 0.995000 ;
      RECT 0.615000  0.995000 1.215000 1.325000 ;
      RECT 0.615000  1.325000 0.785000 2.065000 ;
      RECT 1.035000  0.085000 1.285000 0.585000 ;
      RECT 1.035000  1.575000 1.625000 1.745000 ;
      RECT 1.035000  1.745000 1.365000 2.450000 ;
      RECT 1.455000  0.655000 3.265000 0.825000 ;
      RECT 1.455000  0.825000 1.625000 1.575000 ;
      RECT 1.615000  0.305000 1.785000 0.655000 ;
      RECT 1.985000  0.085000 2.315000 0.485000 ;
      RECT 2.485000  0.305000 2.655000 0.655000 ;
      RECT 2.875000  0.085000 3.255000 0.485000 ;
      RECT 2.920000  1.795000 3.170000 2.635000 ;
      RECT 3.095000  0.825000 3.265000 1.075000 ;
      RECT 3.095000  1.075000 4.555000 1.245000 ;
      RECT 3.815000  1.795000 4.065000 2.635000 ;
      RECT 3.855000  0.085000 4.025000 0.555000 ;
      RECT 4.655000  1.795000 4.905000 2.635000 ;
      RECT 4.695000  0.085000 4.865000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__or4b_4
MACRO sky130_fd_sc_hd__or4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.430000 0.995000 2.810000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 2.125000 2.660000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 0.995000 2.260000 1.615000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.755000 0.425000 1.325000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.320000 0.415000 3.595000 0.760000 ;
        RECT 3.320000 1.495000 3.595000 2.465000 ;
        RECT 3.425000 0.760000 3.595000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.085000 0.425000 0.585000 ;
      RECT 0.085000  1.560000 0.425000 2.635000 ;
      RECT 0.595000  0.305000 0.840000 0.995000 ;
      RECT 0.595000  0.995000 1.250000 1.325000 ;
      RECT 0.595000  1.325000 0.835000 1.920000 ;
      RECT 1.030000  1.495000 1.350000 1.785000 ;
      RECT 1.030000  1.785000 2.660000 1.955000 ;
      RECT 1.035000  0.085000 1.365000 0.585000 ;
      RECT 1.565000  0.305000 1.735000 0.655000 ;
      RECT 1.565000  0.655000 3.150000 0.825000 ;
      RECT 1.910000  0.085000 2.240000 0.485000 ;
      RECT 2.410000  0.305000 2.580000 0.655000 ;
      RECT 2.490000  1.495000 3.150000 1.665000 ;
      RECT 2.490000  1.665000 2.660000 1.785000 ;
      RECT 2.750000  0.085000 3.130000 0.485000 ;
      RECT 2.830000  1.835000 3.110000 2.635000 ;
      RECT 2.980000  0.825000 3.150000 0.995000 ;
      RECT 2.980000  0.995000 3.255000 1.325000 ;
      RECT 2.980000  1.325000 3.150000 1.495000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__or4b_1
MACRO sky130_fd_sc_hd__or4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.755000 1.075000 2.320000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 2.125000 2.670000 2.415000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.550000 1.075000 3.550000 1.275000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.435000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935000 0.675000 1.250000 0.680000 ;
        RECT 0.935000 0.680000 1.245000 0.790000 ;
        RECT 0.935000 0.790000 1.105000 1.495000 ;
        RECT 0.935000 1.495000 1.250000 1.825000 ;
        RECT 0.970000 0.260000 1.250000 0.675000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.325000 0.350000 0.735000 ;
      RECT 0.085000  0.735000 0.765000 0.905000 ;
      RECT 0.085000  1.605000 0.765000 1.890000 ;
      RECT 0.510000  1.890000 0.765000 1.995000 ;
      RECT 0.510000  1.995000 1.715000 2.165000 ;
      RECT 0.515000  2.335000 0.845000 2.635000 ;
      RECT 0.595000  0.905000 0.765000 1.605000 ;
      RECT 0.630000  0.085000 0.800000 0.565000 ;
      RECT 1.290000  0.995000 1.585000 1.325000 ;
      RECT 1.415000  0.735000 3.055000 0.905000 ;
      RECT 1.415000  0.905000 1.585000 0.995000 ;
      RECT 1.415000  1.325000 1.585000 1.355000 ;
      RECT 1.415000  1.355000 1.600000 1.370000 ;
      RECT 1.415000  1.370000 1.610000 1.380000 ;
      RECT 1.415000  1.380000 1.620000 1.390000 ;
      RECT 1.415000  1.390000 1.625000 1.400000 ;
      RECT 1.415000  1.400000 1.630000 1.410000 ;
      RECT 1.415000  1.410000 1.645000 1.420000 ;
      RECT 1.415000  1.420000 1.655000 1.425000 ;
      RECT 1.415000  1.425000 1.665000 1.445000 ;
      RECT 1.415000  1.445000 3.560000 1.450000 ;
      RECT 1.420000  1.450000 3.560000 1.615000 ;
      RECT 1.435000  0.085000 1.815000 0.485000 ;
      RECT 1.440000  1.785000 3.030000 1.955000 ;
      RECT 1.440000  1.955000 1.715000 1.995000 ;
      RECT 1.480000  2.335000 1.815000 2.635000 ;
      RECT 1.985000  0.305000 2.155000 0.735000 ;
      RECT 2.385000  0.085000 2.715000 0.485000 ;
      RECT 2.860000  1.955000 3.030000 2.215000 ;
      RECT 2.860000  2.215000 3.345000 2.385000 ;
      RECT 2.885000  0.305000 3.055000 0.735000 ;
      RECT 3.225000  0.085000 3.555000 0.585000 ;
      RECT 3.225000  1.615000 3.560000 1.815000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__or4b_2
MACRO sky130_fd_sc_hd__a21bo_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21bo_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.750000 0.995000 2.175000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.370000 0.995000 2.630000 1.615000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.325000 0.335000 1.665000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.300000 0.265000 3.580000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.105000  1.845000 0.855000 2.045000 ;
      RECT 0.105000  2.045000 0.345000 2.435000 ;
      RECT 0.515000  0.265000 0.745000 1.165000 ;
      RECT 0.515000  1.165000 0.855000 1.845000 ;
      RECT 0.515000  2.225000 0.865000 2.635000 ;
      RECT 0.945000  0.085000 1.190000 0.865000 ;
      RECT 1.035000  1.045000 1.580000 1.345000 ;
      RECT 1.035000  1.345000 1.365000 2.455000 ;
      RECT 1.360000  0.265000 1.790000 0.625000 ;
      RECT 1.360000  0.625000 3.100000 0.815000 ;
      RECT 1.360000  0.815000 1.580000 1.045000 ;
      RECT 1.535000  1.785000 2.560000 1.985000 ;
      RECT 1.535000  1.985000 1.715000 2.455000 ;
      RECT 1.885000  2.155000 2.215000 2.635000 ;
      RECT 2.370000  0.085000 3.100000 0.455000 ;
      RECT 2.390000  1.985000 2.560000 2.455000 ;
      RECT 2.825000  1.495000 3.110000 2.635000 ;
      RECT 2.840000  0.815000 3.100000 1.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a21bo_1
MACRO sky130_fd_sc_hd__a21bo_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21bo_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685000 0.995000 3.100000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.270000 0.995000 3.560000 1.615000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 1.035000 1.525000 1.325000 ;
        RECT 1.330000 0.995000 1.525000 1.035000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.715000 0.850000 0.885000 ;
        RECT 0.150000 0.885000 0.380000 1.835000 ;
        RECT 0.150000 1.835000 0.850000 2.005000 ;
        RECT 0.520000 0.315000 0.850000 0.715000 ;
        RECT 0.595000 2.005000 0.850000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.090000  0.085000 0.345000 0.545000 ;
      RECT 0.090000  2.255000 0.425000 2.635000 ;
      RECT 0.570000  1.075000 0.900000 1.495000 ;
      RECT 0.570000  1.495000 1.285000 1.665000 ;
      RECT 1.020000  0.085000 1.220000 0.865000 ;
      RECT 1.040000  2.275000 1.370000 2.635000 ;
      RECT 1.115000  1.665000 1.285000 1.895000 ;
      RECT 1.115000  1.895000 2.225000 2.105000 ;
      RECT 1.455000  0.655000 1.865000 0.825000 ;
      RECT 1.455000  1.555000 1.865000 1.725000 ;
      RECT 1.695000  0.825000 1.865000 0.995000 ;
      RECT 1.695000  0.995000 2.175000 1.325000 ;
      RECT 1.695000  1.325000 1.865000 1.555000 ;
      RECT 1.975000  0.085000 2.305000 0.465000 ;
      RECT 1.975000  2.105000 2.225000 2.465000 ;
      RECT 2.055000  1.505000 2.515000 1.675000 ;
      RECT 2.055000  1.675000 2.225000 1.895000 ;
      RECT 2.345000  0.635000 2.740000 0.825000 ;
      RECT 2.345000  0.825000 2.515000 1.505000 ;
      RECT 2.395000  1.845000 3.565000 2.015000 ;
      RECT 2.395000  2.015000 2.725000 2.465000 ;
      RECT 2.895000  2.185000 3.065000 2.635000 ;
      RECT 3.235000  0.085000 3.565000 0.825000 ;
      RECT 3.235000  2.015000 3.565000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__a21bo_2
MACRO sky130_fd_sc_hd__a21bo_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21bo_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.590000 1.010000 4.955000 1.360000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.025000 1.010000 4.420000 1.275000 ;
        RECT 4.245000 1.275000 4.420000 1.595000 ;
        RECT 4.245000 1.595000 5.390000 1.765000 ;
        RECT 5.220000 1.055000 5.700000 1.290000 ;
        RECT 5.220000 1.290000 5.390000 1.595000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.500000 1.010000 0.830000 1.625000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.615000 2.340000 0.785000 ;
        RECT 1.000000 0.785000 1.235000 1.595000 ;
        RECT 1.000000 1.595000 2.410000 1.765000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.105000  0.255000 0.540000 0.840000 ;
      RECT 0.105000  0.840000 0.330000 1.795000 ;
      RECT 0.105000  1.795000 0.565000 1.935000 ;
      RECT 0.105000  1.935000 2.870000 2.105000 ;
      RECT 0.105000  2.105000 0.550000 2.465000 ;
      RECT 0.710000  0.085000 1.050000 0.445000 ;
      RECT 0.720000  2.275000 1.050000 2.635000 ;
      RECT 1.405000  0.995000 2.810000 1.185000 ;
      RECT 1.405000  1.185000 2.530000 1.325000 ;
      RECT 1.580000  0.085000 1.910000 0.445000 ;
      RECT 1.580000  2.275000 1.910000 2.635000 ;
      RECT 2.435000  2.275000 2.770000 2.635000 ;
      RECT 2.515000  0.085000 3.285000 0.445000 ;
      RECT 2.640000  0.615000 3.645000 0.670000 ;
      RECT 2.640000  0.670000 4.965000 0.785000 ;
      RECT 2.640000  0.785000 3.010000 0.800000 ;
      RECT 2.640000  0.800000 2.810000 0.995000 ;
      RECT 2.700000  1.355000 3.305000 1.525000 ;
      RECT 2.700000  1.525000 2.870000 1.935000 ;
      RECT 2.995000  0.995000 3.305000 1.355000 ;
      RECT 3.055000  1.695000 3.225000 2.210000 ;
      RECT 3.055000  2.210000 4.065000 2.380000 ;
      RECT 3.475000  0.255000 3.645000 0.615000 ;
      RECT 3.475000  0.785000 4.965000 0.840000 ;
      RECT 3.475000  0.840000 3.645000 1.805000 ;
      RECT 3.855000  0.085000 4.185000 0.445000 ;
      RECT 3.885000  1.445000 4.065000 1.935000 ;
      RECT 3.885000  1.935000 5.825000 2.105000 ;
      RECT 3.885000  2.105000 4.065000 2.210000 ;
      RECT 4.235000  2.275000 4.565000 2.635000 ;
      RECT 4.685000  0.405000 4.965000 0.670000 ;
      RECT 5.075000  2.275000 5.405000 2.635000 ;
      RECT 5.545000  0.085000 5.825000 0.885000 ;
      RECT 5.570000  1.460000 5.825000 1.935000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
END sky130_fd_sc_hd__a21bo_4
MACRO sky130_fd_sc_hd__nand2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.440000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155000 1.075000 4.940000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 0.635000 2.640000 0.905000 ;
        RECT 1.455000 1.445000 4.320000 1.665000 ;
        RECT 1.455000 1.665000 1.785000 2.465000 ;
        RECT 2.295000 1.665000 2.640000 2.465000 ;
        RECT 2.375000 0.905000 2.640000 1.445000 ;
        RECT 3.150000 1.665000 3.480000 2.465000 ;
        RECT 3.990000 1.665000 4.320000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.060000 0.085000 ;
      RECT 0.000000  2.635000 5.060000 2.805000 ;
      RECT 0.090000  0.255000 0.425000 0.715000 ;
      RECT 0.090000  0.715000 0.780000 0.905000 ;
      RECT 0.090000  1.445000 0.780000 1.665000 ;
      RECT 0.090000  1.665000 0.425000 2.465000 ;
      RECT 0.595000  0.085000 0.790000 0.545000 ;
      RECT 0.595000  1.835000 1.285000 2.635000 ;
      RECT 0.610000  0.905000 0.780000 1.075000 ;
      RECT 0.610000  1.075000 2.205000 1.275000 ;
      RECT 0.610000  1.275000 0.780000 1.445000 ;
      RECT 0.970000  1.445000 1.285000 1.835000 ;
      RECT 1.035000  0.255000 3.060000 0.465000 ;
      RECT 1.035000  0.465000 1.285000 0.905000 ;
      RECT 1.955000  1.835000 2.125000 2.635000 ;
      RECT 2.810000  0.465000 3.060000 0.715000 ;
      RECT 2.810000  0.715000 4.850000 0.905000 ;
      RECT 2.810000  1.835000 2.980000 2.635000 ;
      RECT 3.230000  0.085000 3.400000 0.545000 ;
      RECT 3.570000  0.255000 3.900000 0.715000 ;
      RECT 3.650000  1.835000 3.820000 2.635000 ;
      RECT 4.070000  0.085000 4.310000 0.545000 ;
      RECT 4.520000  0.255000 4.850000 0.715000 ;
      RECT 4.520000  1.495000 4.850000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2b_4
MACRO sky130_fd_sc_hd__nand2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.440000 1.315000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.075000 1.085000 1.315000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 1.835000 2.170000 2.005000 ;
        RECT 1.000000 2.005000 1.330000 2.465000 ;
        RECT 1.420000 0.255000 2.170000 0.545000 ;
        RECT 1.800000 0.545000 2.170000 1.835000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.090000  0.525000 0.360000 0.735000 ;
      RECT 0.090000  0.735000 1.425000 0.905000 ;
      RECT 0.090000  1.495000 1.425000 1.665000 ;
      RECT 0.090000  1.665000 0.370000 1.825000 ;
      RECT 0.580000  0.085000 0.910000 0.545000 ;
      RECT 0.580000  1.835000 0.830000 2.635000 ;
      RECT 1.255000  0.905000 1.425000 1.075000 ;
      RECT 1.255000  1.075000 1.630000 1.325000 ;
      RECT 1.255000  1.325000 1.425000 1.495000 ;
      RECT 1.500000  2.175000 1.715000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2b_1
MACRO sky130_fd_sc_hd__nand2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 0.995000 0.800000 1.325000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.075000 3.135000 1.275000 ;
        RECT 1.990000 1.275000 2.180000 1.655000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.775500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.835000 2.635000 2.005000 ;
        RECT 1.035000 2.005000 1.365000 2.465000 ;
        RECT 1.525000 0.635000 1.855000 0.805000 ;
        RECT 1.530000 0.805000 1.855000 0.905000 ;
        RECT 1.530000 0.905000 1.810000 1.835000 ;
        RECT 2.280000 2.005000 2.635000 2.465000 ;
        RECT 2.360000 1.495000 2.635000 1.835000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.110000  0.510000 0.345000 0.840000 ;
      RECT 0.110000  0.840000 0.280000 1.495000 ;
      RECT 0.110000  1.495000 1.360000 1.665000 ;
      RECT 0.110000  1.665000 0.410000 1.860000 ;
      RECT 0.515000  0.085000 0.845000 0.825000 ;
      RECT 0.580000  1.835000 0.835000 2.635000 ;
      RECT 1.030000  1.075000 1.360000 1.495000 ;
      RECT 1.080000  0.255000 2.275000 0.465000 ;
      RECT 1.080000  0.465000 1.355000 0.905000 ;
      RECT 1.535000  2.175000 2.110000 2.635000 ;
      RECT 2.025000  0.465000 2.275000 0.695000 ;
      RECT 2.025000  0.695000 3.135000 0.905000 ;
      RECT 2.445000  0.085000 2.615000 0.525000 ;
      RECT 2.785000  0.255000 3.135000 0.695000 ;
      RECT 2.805000  1.495000 3.135000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__nand2b_2
MACRO sky130_fd_sc_hd__nor3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 0.995000 1.815000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.995000 1.305000 1.615000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.995000 2.335000 1.615000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  0.716500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.605000 0.655000 ;
        RECT 0.085000 0.655000 1.445000 0.825000 ;
        RECT 0.085000 0.825000 0.255000 1.445000 ;
        RECT 0.085000 1.445000 0.545000 2.455000 ;
        RECT 1.275000 0.310000 1.445000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.950000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.425000  1.075000 0.885000 1.245000 ;
      RECT 0.715000  1.245000 0.885000 1.785000 ;
      RECT 0.715000  1.785000 2.675000 1.955000 ;
      RECT 0.775000  0.085000 1.105000 0.485000 ;
      RECT 1.615000  0.085000 1.945000 0.825000 ;
      RECT 1.615000  2.125000 1.945000 2.635000 ;
      RECT 2.180000  0.405000 2.350000 0.655000 ;
      RECT 2.180000  0.655000 2.675000 0.825000 ;
      RECT 2.505000  0.825000 2.675000 1.785000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
END sky130_fd_sc_hd__nor3b_1
MACRO sky130_fd_sc_hd__nor3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.075000 2.690000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 1.075000 4.300000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.445000 1.285000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 0.255000 1.285000 0.725000 ;
        RECT 0.955000 0.725000 6.760000 0.905000 ;
        RECT 1.795000 0.255000 2.125000 0.725000 ;
        RECT 3.155000 0.255000 3.485000 0.725000 ;
        RECT 3.995000 0.255000 4.325000 0.725000 ;
        RECT 4.835000 0.255000 5.165000 0.725000 ;
        RECT 4.875000 1.455000 6.760000 1.625000 ;
        RECT 4.875000 1.625000 5.125000 2.125000 ;
        RECT 5.675000 0.255000 6.005000 0.725000 ;
        RECT 5.715000 1.625000 5.965000 2.125000 ;
        RECT 6.420000 0.905000 6.760000 1.455000 ;
        RECT 6.515000 0.315000 6.760000 0.725000 ;
        RECT 6.555000 1.625000 6.760000 2.415000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.090000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.900000 0.085000 ;
      RECT 0.000000  2.635000 6.900000 2.805000 ;
      RECT 0.110000  0.255000 0.445000 0.735000 ;
      RECT 0.110000  0.735000 0.785000 0.905000 ;
      RECT 0.110000  1.455000 4.705000 1.625000 ;
      RECT 0.110000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.615000  0.085000 0.785000 0.555000 ;
      RECT 0.615000  0.905000 0.785000 1.455000 ;
      RECT 0.995000  1.795000 4.285000 1.965000 ;
      RECT 0.995000  1.965000 1.245000 2.465000 ;
      RECT 1.415000  2.135000 1.665000 2.635000 ;
      RECT 1.455000  0.085000 1.625000 0.555000 ;
      RECT 1.835000  1.965000 2.085000 2.465000 ;
      RECT 2.255000  2.135000 2.505000 2.635000 ;
      RECT 2.295000  0.085000 2.985000 0.555000 ;
      RECT 2.775000  2.135000 3.025000 2.295000 ;
      RECT 2.775000  2.295000 6.385000 2.465000 ;
      RECT 3.195000  1.965000 3.445000 2.125000 ;
      RECT 3.615000  2.135000 3.865000 2.295000 ;
      RECT 3.655000  0.085000 3.825000 0.555000 ;
      RECT 4.035000  1.965000 4.285000 2.125000 ;
      RECT 4.455000  1.795000 4.705000 2.295000 ;
      RECT 4.495000  0.085000 4.665000 0.555000 ;
      RECT 4.535000  1.075000 6.125000 1.285000 ;
      RECT 4.535000  1.285000 4.705000 1.455000 ;
      RECT 5.295000  1.795000 5.545000 2.295000 ;
      RECT 5.335000  0.085000 5.505000 0.555000 ;
      RECT 6.135000  1.795000 6.385000 2.295000 ;
      RECT 6.175000  0.085000 6.345000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
  END
END sky130_fd_sc_hd__nor3b_4
MACRO sky130_fd_sc_hd__nor3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.965000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135000 1.075000 2.640000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.030000 1.075000 4.515000 1.285000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 3.105000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.775000 0.255000 3.105000 0.725000 ;
        RECT 2.815000 0.905000 3.065000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 2.085000 1.625000 ;
      RECT 0.090000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.995000  1.625000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.795000 1.665000 2.295000 ;
      RECT 1.415000  2.295000 3.480000 2.465000 ;
      RECT 1.835000  1.625000 2.085000 2.125000 ;
      RECT 1.875000  0.085000 2.605000 0.555000 ;
      RECT 2.375000  1.455000 2.645000 2.295000 ;
      RECT 3.235000  1.075000 3.860000 1.285000 ;
      RECT 3.235000  1.455000 3.480000 2.295000 ;
      RECT 3.275000  0.085000 3.480000 0.895000 ;
      RECT 3.690000  0.380000 4.045000 0.905000 ;
      RECT 3.690000  0.905000 3.860000 1.075000 ;
      RECT 3.690000  1.285000 3.860000 1.455000 ;
      RECT 3.690000  1.455000 4.045000 1.870000 ;
      RECT 4.215000  0.085000 4.505000 0.825000 ;
      RECT 4.215000  1.540000 4.465000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__nor3b_2
MACRO sky130_fd_sc_hd__o22ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 1.075000 4.165000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.075000 3.225000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.200000 1.075000 0.985000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.155000 1.075000 1.925000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.645000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 2.340000 0.905000 ;
        RECT 1.375000 0.645000 1.705000 0.725000 ;
        RECT 1.415000 1.445000 3.065000 1.625000 ;
        RECT 1.415000 1.625000 1.665000 2.125000 ;
        RECT 2.095000 0.905000 2.340000 1.445000 ;
        RECT 2.815000 1.625000 3.065000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.305000 2.680000 0.475000 ;
      RECT 0.090000  0.475000 0.365000 0.905000 ;
      RECT 0.150000  1.455000 1.245000 1.625000 ;
      RECT 0.150000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.995000  1.625000 1.245000 2.295000 ;
      RECT 0.995000  2.295000 2.085000 2.465000 ;
      RECT 1.835000  1.795000 2.085000 2.295000 ;
      RECT 2.395000  1.795000 2.645000 2.295000 ;
      RECT 2.395000  2.295000 3.485000 2.465000 ;
      RECT 2.510000  0.475000 2.680000 0.725000 ;
      RECT 2.510000  0.725000 4.365000 0.905000 ;
      RECT 2.855000  0.085000 3.025000 0.555000 ;
      RECT 3.195000  0.255000 3.525000 0.725000 ;
      RECT 3.235000  1.455000 4.330000 1.625000 ;
      RECT 3.235000  1.625000 3.485000 2.295000 ;
      RECT 3.655000  1.795000 3.905000 2.635000 ;
      RECT 3.695000  0.085000 3.865000 0.555000 ;
      RECT 4.035000  0.255000 4.365000 0.725000 ;
      RECT 4.075000  1.625000 4.330000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__o22ai_2
MACRO sky130_fd_sc_hd__o22ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.755000 1.075000 2.215000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.220000 1.075000 1.585000 1.245000 ;
        RECT 1.405000 1.245000 1.585000 1.445000 ;
        RECT 1.405000 1.445000 1.725000 1.615000 ;
        RECT 1.525000 1.615000 1.725000 2.405000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.665000 0.325000 1.990000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 0.995000 1.005000 1.415000 ;
        RECT 0.835000 1.415000 1.235000 1.665000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.650250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495000 0.645000 0.845000 0.825000 ;
        RECT 0.495000 0.825000 0.665000 1.835000 ;
        RECT 0.495000 1.835000 1.335000 2.045000 ;
        RECT 0.835000 2.045000 1.335000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.295000 1.345000 0.475000 ;
      RECT 0.135000  2.175000 0.345000 2.635000 ;
      RECT 1.015000  0.475000 1.345000 0.695000 ;
      RECT 1.015000  0.695000 2.215000 0.825000 ;
      RECT 1.185000  0.825000 2.215000 0.865000 ;
      RECT 1.535000  0.085000 1.705000 0.525000 ;
      RECT 1.875000  0.280000 2.215000 0.695000 ;
      RECT 1.895000  1.455000 2.215000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__o22ai_1
MACRO sky130_fd_sc_hd__o22ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 1.415000 1.275000 ;
        RECT 1.150000 1.275000 1.415000 1.445000 ;
        RECT 1.150000 1.445000 3.575000 1.615000 ;
        RECT 3.275000 1.075000 3.605000 1.245000 ;
        RECT 3.275000 1.245000 3.575000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.685000 1.075000 3.095000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.295000 0.995000 4.940000 1.445000 ;
        RECT 4.295000 1.445000 6.935000 1.615000 ;
        RECT 6.715000 0.995000 6.935000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.110000 1.075000 6.460000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845000 1.785000 3.915000 1.955000 ;
        RECT 1.845000 1.955000 2.095000 2.125000 ;
        RECT 2.685000 1.955000 2.935000 2.125000 ;
        RECT 3.745000 1.445000 4.125000 1.615000 ;
        RECT 3.745000 1.615000 3.915000 1.785000 ;
        RECT 3.955000 0.645000 7.275000 0.820000 ;
        RECT 3.955000 0.820000 4.125000 1.445000 ;
        RECT 5.255000 1.785000 7.275000 1.955000 ;
        RECT 5.255000 1.955000 5.505000 2.125000 ;
        RECT 6.095000 1.955000 6.345000 2.125000 ;
        RECT 7.105000 0.820000 7.275000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.125000  0.255000 0.455000 0.725000 ;
      RECT 0.125000  0.725000 1.295000 0.735000 ;
      RECT 0.125000  0.735000 3.785000 0.905000 ;
      RECT 0.165000  1.445000 0.415000 2.635000 ;
      RECT 0.585000  1.445000 0.835000 1.785000 ;
      RECT 0.585000  1.785000 1.675000 1.955000 ;
      RECT 0.585000  1.955000 0.835000 2.465000 ;
      RECT 0.625000  0.085000 0.795000 0.555000 ;
      RECT 0.965000  0.255000 1.295000 0.725000 ;
      RECT 1.005000  2.125000 1.255000 2.635000 ;
      RECT 1.425000  1.955000 1.675000 2.295000 ;
      RECT 1.425000  2.295000 3.395000 2.465000 ;
      RECT 1.465000  0.085000 1.635000 0.555000 ;
      RECT 1.805000  0.255000 2.135000 0.725000 ;
      RECT 1.805000  0.725000 2.975000 0.735000 ;
      RECT 2.265000  2.125000 2.515000 2.295000 ;
      RECT 2.305000  0.085000 2.475000 0.555000 ;
      RECT 2.645000  0.255000 2.975000 0.725000 ;
      RECT 3.105000  2.125000 3.395000 2.295000 ;
      RECT 3.145000  0.085000 3.315000 0.555000 ;
      RECT 3.485000  0.255000 7.245000 0.475000 ;
      RECT 3.485000  0.475000 3.785000 0.735000 ;
      RECT 3.565000  2.125000 3.785000 2.635000 ;
      RECT 3.955000  2.125000 4.255000 2.465000 ;
      RECT 4.085000  1.785000 5.085000 1.955000 ;
      RECT 4.085000  1.955000 4.255000 2.125000 ;
      RECT 4.425000  2.125000 4.665000 2.635000 ;
      RECT 4.835000  1.955000 5.085000 2.295000 ;
      RECT 4.835000  2.295000 6.765000 2.465000 ;
      RECT 5.675000  2.125000 5.925000 2.295000 ;
      RECT 6.515000  2.135000 6.765000 2.295000 ;
      RECT 6.935000  2.125000 7.215000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__o22ai_4
MACRO sky130_fd_sc_hd__o2bb2ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095000 1.075000 3.505000 1.285000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 1.825000 1.285000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.045000 1.075000 10.005000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465000 1.075000 7.875000 1.285000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.415000 0.645000 6.155000 0.905000 ;
        RECT 4.425000 1.455000 7.715000 1.625000 ;
        RECT 4.425000 1.625000 4.675000 2.465000 ;
        RECT 5.265000 1.625000 5.515000 2.465000 ;
        RECT 5.875000 0.905000 6.155000 1.455000 ;
        RECT 6.625000 1.625000 6.875000 2.125000 ;
        RECT 7.465000 1.625000 7.715000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.135000 -0.085000 0.305000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.310000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.120000 0.085000 ;
      RECT 0.000000  2.635000 10.120000 2.805000 ;
      RECT 0.085000  0.645000  1.705000 0.905000 ;
      RECT 0.085000  0.905000  0.255000 1.455000 ;
      RECT 0.085000  1.455000  3.915000 1.625000 ;
      RECT 0.100000  0.255000  2.125000 0.475000 ;
      RECT 0.155000  1.795000  0.405000 2.635000 ;
      RECT 0.575000  1.625000  0.825000 2.465000 ;
      RECT 0.995000  1.795000  1.245000 2.635000 ;
      RECT 1.415000  1.625000  1.665000 2.465000 ;
      RECT 1.835000  1.795000  2.085000 2.635000 ;
      RECT 1.875000  0.475000  2.125000 0.725000 ;
      RECT 1.875000  0.725000  3.805000 0.905000 ;
      RECT 2.255000  1.625000  2.505000 2.465000 ;
      RECT 2.295000  0.085000  2.465000 0.555000 ;
      RECT 2.635000  0.255000  2.965000 0.725000 ;
      RECT 2.675000  1.795000  2.925000 2.635000 ;
      RECT 3.095000  1.625000  3.345000 2.465000 ;
      RECT 3.135000  0.085000  3.305000 0.555000 ;
      RECT 3.475000  0.255000  3.805000 0.725000 ;
      RECT 3.515000  1.795000  4.255000 2.635000 ;
      RECT 3.745000  1.075000  5.705000 1.285000 ;
      RECT 3.745000  1.285000  3.915000 1.455000 ;
      RECT 4.060000  0.255000  6.495000 0.475000 ;
      RECT 4.060000  0.475000  4.245000 0.835000 ;
      RECT 4.845000  1.795000  5.095000 2.635000 ;
      RECT 5.685000  1.795000  5.935000 2.635000 ;
      RECT 6.175000  1.795000  6.455000 2.295000 ;
      RECT 6.175000  2.295000  8.135000 2.465000 ;
      RECT 6.325000  0.475000  6.495000 0.735000 ;
      RECT 6.325000  0.735000  9.855000 0.905000 ;
      RECT 6.665000  0.085000  6.835000 0.555000 ;
      RECT 7.005000  0.255000  7.335000 0.725000 ;
      RECT 7.005000  0.725000  9.855000 0.735000 ;
      RECT 7.045000  1.795000  7.295000 2.295000 ;
      RECT 7.505000  0.085000  7.675000 0.555000 ;
      RECT 7.845000  0.255000  8.175000 0.725000 ;
      RECT 7.885000  1.455000  9.875000 1.625000 ;
      RECT 7.885000  1.625000  8.135000 2.295000 ;
      RECT 8.305000  1.795000  8.555000 2.635000 ;
      RECT 8.345000  0.085000  8.515000 0.555000 ;
      RECT 8.685000  0.255000  9.015000 0.725000 ;
      RECT 8.725000  1.625000  8.975000 2.465000 ;
      RECT 9.145000  1.795000  9.395000 2.635000 ;
      RECT 9.185000  0.085000  9.355000 0.555000 ;
      RECT 9.525000  0.255000  9.855000 0.725000 ;
      RECT 9.565000  1.625000  9.875000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
      RECT 9.805000 -0.085000 9.975000 0.085000 ;
      RECT 9.805000  2.635000 9.975000 2.805000 ;
  END
END sky130_fd_sc_hd__o2bb2ai_4
MACRO sky130_fd_sc_hd__o2bb2ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.625000 1.445000 ;
        RECT 0.090000 1.445000 1.945000 1.615000 ;
        RECT 1.615000 1.075000 1.945000 1.445000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.795000 1.075000 1.400000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.410000 1.075000 3.740000 1.445000 ;
        RECT 3.410000 1.445000 5.435000 1.615000 ;
        RECT 4.730000 1.075000 5.435000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.960000 1.075000 4.500000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.745000 0.645000 3.075000 1.075000 ;
        RECT 2.745000 1.075000 3.215000 1.785000 ;
        RECT 2.745000 1.785000 4.330000 1.955000 ;
        RECT 2.745000 1.955000 3.035000 2.465000 ;
        RECT 4.080000 1.955000 4.330000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.150000  1.795000 0.400000 2.635000 ;
      RECT 0.195000  0.085000 0.365000 0.895000 ;
      RECT 0.535000  0.305000 1.705000 0.475000 ;
      RECT 0.535000  0.475000 0.785000 0.895000 ;
      RECT 0.575000  1.785000 2.285000 1.965000 ;
      RECT 0.575000  1.965000 0.825000 2.465000 ;
      RECT 0.955000  0.645000 1.285000 0.725000 ;
      RECT 0.955000  0.725000 2.285000 0.905000 ;
      RECT 0.995000  2.135000 1.245000 2.635000 ;
      RECT 1.415000  1.965000 1.665000 2.125000 ;
      RECT 1.835000  2.135000 2.575000 2.635000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.115000  0.905000 2.285000 0.995000 ;
      RECT 2.115000  0.995000 2.575000 1.325000 ;
      RECT 2.115000  1.325000 2.285000 1.785000 ;
      RECT 2.325000  0.255000 3.530000 0.475000 ;
      RECT 2.325000  0.475000 2.575000 0.555000 ;
      RECT 3.205000  2.125000 3.490000 2.635000 ;
      RECT 3.245000  0.475000 3.530000 0.735000 ;
      RECT 3.245000  0.735000 5.210000 0.905000 ;
      RECT 3.660000  2.125000 3.910000 2.295000 ;
      RECT 3.660000  2.295000 4.750000 2.465000 ;
      RECT 3.700000  0.085000 3.870000 0.555000 ;
      RECT 4.040000  0.255000 4.370000 0.725000 ;
      RECT 4.040000  0.725000 5.210000 0.735000 ;
      RECT 4.500000  1.785000 4.750000 2.295000 ;
      RECT 4.540000  0.085000 4.710000 0.555000 ;
      RECT 4.880000  0.255000 5.210000 0.725000 ;
      RECT 4.965000  1.795000 5.170000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__o2bb2ai_2
MACRO sky130_fd_sc_hd__o2bb2ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.435000 1.285000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.280000 0.825000 0.995000 ;
        RECT 0.605000 0.995000 1.000000 1.325000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 1.075000 3.135000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.030000 1.075000 2.615000 1.325000 ;
        RECT 2.445000 1.325000 2.615000 2.425000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.560000 0.430000 1.810000 0.790000 ;
        RECT 1.640000 0.790000 1.810000 1.495000 ;
        RECT 1.640000 1.495000 2.270000 1.665000 ;
        RECT 1.940000 1.665000 2.270000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.090000  0.085000 0.425000 0.815000 ;
      RECT 0.150000  1.455000 0.400000 2.635000 ;
      RECT 0.570000  1.495000 1.340000 1.665000 ;
      RECT 0.570000  1.665000 0.820000 2.465000 ;
      RECT 0.990000  1.835000 1.770000 2.635000 ;
      RECT 1.000000  0.280000 1.340000 0.825000 ;
      RECT 1.170000  0.825000 1.340000 0.995000 ;
      RECT 1.170000  0.995000 1.470000 1.325000 ;
      RECT 1.170000  1.325000 1.340000 1.495000 ;
      RECT 1.980000  0.425000 2.270000 0.725000 ;
      RECT 1.980000  0.725000 3.110000 0.905000 ;
      RECT 2.440000  0.085000 2.610000 0.555000 ;
      RECT 2.780000  0.275000 3.110000 0.725000 ;
      RECT 2.820000  1.455000 3.070000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__o2bb2ai_1
MACRO sky130_fd_sc_hd__sdfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 1.355000 2.775000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.180000 0.305000 9.530000 0.725000 ;
        RECT 9.180000 0.725000 9.560000 0.790000 ;
        RECT 9.180000 0.790000 9.610000 0.825000 ;
        RECT 9.200000 1.505000 9.610000 1.540000 ;
        RECT 9.200000 1.540000 9.530000 2.465000 ;
        RECT 9.355000 1.430000 9.610000 1.505000 ;
        RECT 9.390000 0.825000 9.610000 1.430000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685000 0.265000 10.940000 0.795000 ;
        RECT 10.685000 1.445000 10.940000 2.325000 ;
        RECT 10.730000 0.795000 10.940000 1.445000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515000 1.055000 3.995000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.760000 0.750000 3.235000 0.785000 ;
        RECT 1.760000 0.785000 2.010000 0.810000 ;
        RECT 1.760000 0.810000 1.990000 0.820000 ;
        RECT 1.760000 0.820000 1.975000 0.835000 ;
        RECT 1.760000 0.835000 1.970000 0.840000 ;
        RECT 1.760000 0.840000 1.965000 0.850000 ;
        RECT 1.760000 0.850000 1.960000 0.855000 ;
        RECT 1.760000 0.855000 1.955000 0.860000 ;
        RECT 1.760000 0.860000 1.950000 0.870000 ;
        RECT 1.760000 0.870000 1.945000 0.875000 ;
        RECT 1.760000 0.875000 1.940000 0.880000 ;
        RECT 1.760000 0.880000 1.930000 1.685000 ;
        RECT 1.790000 0.735000 3.235000 0.750000 ;
        RECT 1.805000 0.725000 3.235000 0.735000 ;
        RECT 1.820000 0.715000 3.235000 0.725000 ;
        RECT 1.830000 0.705000 3.235000 0.715000 ;
        RECT 1.840000 0.690000 3.235000 0.705000 ;
        RECT 1.860000 0.655000 3.235000 0.690000 ;
        RECT 1.875000 0.615000 3.235000 0.655000 ;
        RECT 2.455000 0.305000 2.630000 0.615000 ;
        RECT 3.065000 0.785000 3.235000 1.115000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 11.230000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  2.635000 11.040000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.810000 0.805000 ;
      RECT  0.175000  1.795000  0.845000 1.965000 ;
      RECT  0.175000  1.965000  0.345000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.515000  2.135000  0.845000 2.635000 ;
      RECT  0.615000  0.805000  0.810000 0.970000 ;
      RECT  0.615000  0.970000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.185000 2.465000 ;
      RECT  1.420000  0.255000  1.705000 0.585000 ;
      RECT  1.420000  0.585000  1.590000 1.860000 ;
      RECT  1.420000  1.860000  3.230000 2.075000 ;
      RECT  1.420000  2.075000  1.705000 2.445000 ;
      RECT  1.875000  2.245000  2.205000 2.635000 ;
      RECT  1.955000  0.085000  2.285000 0.445000 ;
      RECT  2.100000  0.955000  2.445000 1.125000 ;
      RECT  2.100000  1.125000  2.270000 1.860000 ;
      RECT  2.675000  2.245000  3.570000 2.415000 ;
      RECT  2.800000  0.275000  3.575000 0.445000 ;
      RECT  3.060000  1.355000  3.255000 1.685000 ;
      RECT  3.060000  1.685000  3.230000 1.860000 ;
      RECT  3.400000  1.825000  4.335000 1.995000 ;
      RECT  3.400000  1.995000  3.570000 2.245000 ;
      RECT  3.405000  0.445000  3.575000 0.715000 ;
      RECT  3.405000  0.715000  4.335000 0.885000 ;
      RECT  3.740000  2.165000  3.910000 2.635000 ;
      RECT  3.745000  0.085000  3.945000 0.545000 ;
      RECT  4.165000  0.365000  4.515000 0.535000 ;
      RECT  4.165000  0.535000  4.335000 0.715000 ;
      RECT  4.165000  0.885000  4.335000 1.825000 ;
      RECT  4.165000  1.995000  4.335000 2.070000 ;
      RECT  4.165000  2.070000  4.450000 2.440000 ;
      RECT  4.505000  0.705000  5.085000 1.035000 ;
      RECT  4.505000  1.035000  4.745000 1.905000 ;
      RECT  4.645000  2.190000  5.715000 2.360000 ;
      RECT  4.685000  0.365000  5.425000 0.535000 ;
      RECT  4.935000  1.655000  5.375000 2.010000 ;
      RECT  5.255000  0.535000  5.425000 1.315000 ;
      RECT  5.255000  1.315000  6.055000 1.485000 ;
      RECT  5.545000  1.485000  6.055000 1.575000 ;
      RECT  5.545000  1.575000  5.715000 2.190000 ;
      RECT  5.595000  0.765000  6.395000 1.065000 ;
      RECT  5.595000  1.065000  5.765000 1.095000 ;
      RECT  5.675000  0.085000  6.045000 0.585000 ;
      RECT  5.885000  1.245000  6.055000 1.315000 ;
      RECT  5.885000  1.835000  6.055000 2.635000 ;
      RECT  6.225000  0.365000  6.685000 0.535000 ;
      RECT  6.225000  0.535000  6.395000 0.765000 ;
      RECT  6.225000  1.065000  6.395000 2.135000 ;
      RECT  6.225000  2.135000  6.475000 2.465000 ;
      RECT  6.565000  0.705000  7.115000 1.035000 ;
      RECT  6.565000  1.245000  6.755000 1.965000 ;
      RECT  6.700000  2.165000  7.585000 2.335000 ;
      RECT  6.915000  0.365000  7.455000 0.535000 ;
      RECT  6.925000  1.035000  7.115000 1.575000 ;
      RECT  6.925000  1.575000  7.245000 1.905000 ;
      RECT  7.285000  0.535000  7.455000 0.995000 ;
      RECT  7.285000  0.995000  8.315000 1.325000 ;
      RECT  7.285000  1.325000  7.585000 1.405000 ;
      RECT  7.415000  1.405000  7.585000 2.165000 ;
      RECT  7.700000  0.085000  8.070000 0.615000 ;
      RECT  7.755000  1.575000  8.670000 1.905000 ;
      RECT  7.765000  2.135000  8.070000 2.635000 ;
      RECT  8.340000  0.300000  8.670000 0.825000 ;
      RECT  8.380000  1.905000  8.670000 2.455000 ;
      RECT  8.485000  0.825000  8.670000 0.995000 ;
      RECT  8.485000  0.995000  9.220000 1.325000 ;
      RECT  8.485000  1.325000  8.670000 1.575000 ;
      RECT  8.840000  0.085000  9.010000 0.695000 ;
      RECT  8.840000  1.625000  9.010000 2.635000 ;
      RECT  9.700000  0.345000  9.950000 0.620000 ;
      RECT  9.700000  1.685000 10.030000 2.425000 ;
      RECT  9.780000  0.620000  9.950000 0.995000 ;
      RECT  9.780000  0.995000 10.560000 1.325000 ;
      RECT  9.780000  1.325000 10.030000 1.685000 ;
      RECT 10.185000  0.085000 10.515000 0.805000 ;
      RECT 10.210000  1.495000 10.515000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.645000  1.785000  0.815000 1.955000 ;
      RECT  1.015000  0.765000  1.185000 0.935000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  0.765000  4.915000 0.935000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.165000  1.785000  5.335000 1.955000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.575000  1.785000  6.745000 1.955000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  0.765000  6.755000 0.935000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
    LAYER met1 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 6.805000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 0.955000 0.735000 1.245000 0.780000 ;
      RECT 0.955000 0.780000 6.815000 0.920000 ;
      RECT 0.955000 0.920000 1.245000 0.965000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.105000 1.755000 5.395000 1.800000 ;
      RECT 5.105000 1.940000 5.395000 1.985000 ;
      RECT 6.515000 1.755000 6.805000 1.800000 ;
      RECT 6.515000 1.940000 6.805000 1.985000 ;
      RECT 6.525000 0.735000 6.815000 0.780000 ;
      RECT 6.525000 0.920000 6.815000 0.965000 ;
  END
END sky130_fd_sc_hd__sdfxbp_1
MACRO sky130_fd_sc_hd__sdfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.460000 1.355000 2.795000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.255000 0.255000 9.585000 0.790000 ;
        RECT 9.255000 0.790000 9.615000 0.825000 ;
        RECT 9.255000 1.495000 9.615000 1.530000 ;
        RECT 9.255000 1.530000 9.585000 2.430000 ;
        RECT 9.410000 0.825000 9.615000 0.890000 ;
        RECT 9.410000 1.430000 9.615000 1.495000 ;
        RECT 9.445000 0.890000 9.615000 1.430000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.190000 0.265000 11.440000 0.795000 ;
        RECT 11.190000 1.445000 11.440000 2.325000 ;
        RECT 11.235000 0.795000 11.440000 1.445000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.535000 1.035000 4.035000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.615000 3.255000 0.785000 ;
        RECT 1.780000 0.785000 1.950000 1.685000 ;
        RECT 2.475000 0.305000 2.650000 0.615000 ;
        RECT 3.085000 0.785000 3.255000 1.115000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.810000 0.805000 ;
      RECT  0.180000  1.795000  0.845000 1.965000 ;
      RECT  0.180000  1.965000  0.350000 2.465000 ;
      RECT  0.515000  0.085000  0.845000 0.465000 ;
      RECT  0.520000  2.135000  0.850000 2.635000 ;
      RECT  0.615000  0.805000  0.810000 0.970000 ;
      RECT  0.615000  0.970000  0.845000 1.795000 ;
      RECT  1.015000  0.345000  1.245000 0.715000 ;
      RECT  1.020000  0.715000  1.245000 2.465000 ;
      RECT  1.435000  0.275000  1.805000 0.445000 ;
      RECT  1.435000  0.445000  1.605000 1.860000 ;
      RECT  1.435000  1.860000  3.250000 2.075000 ;
      RECT  1.435000  2.075000  1.710000 2.445000 ;
      RECT  1.880000  2.245000  2.210000 2.635000 ;
      RECT  1.975000  0.085000  2.305000 0.445000 ;
      RECT  2.120000  0.955000  2.465000 1.125000 ;
      RECT  2.120000  1.125000  2.290000 1.860000 ;
      RECT  2.695000  2.245000  3.590000 2.415000 ;
      RECT  2.820000  0.275000  3.595000 0.445000 ;
      RECT  3.080000  1.355000  3.275000 1.685000 ;
      RECT  3.080000  1.685000  3.250000 1.860000 ;
      RECT  3.420000  1.825000  4.375000 1.995000 ;
      RECT  3.420000  1.995000  3.590000 2.245000 ;
      RECT  3.425000  0.445000  3.595000 0.695000 ;
      RECT  3.425000  0.695000  4.375000 0.865000 ;
      RECT  3.760000  2.165000  3.930000 2.635000 ;
      RECT  3.765000  0.085000  3.965000 0.525000 ;
      RECT  4.205000  0.365000  4.555000 0.535000 ;
      RECT  4.205000  0.535000  4.375000 0.695000 ;
      RECT  4.205000  0.865000  4.375000 1.825000 ;
      RECT  4.205000  1.995000  4.375000 2.065000 ;
      RECT  4.205000  2.065000  4.485000 2.440000 ;
      RECT  4.545000  0.705000  5.125000 1.035000 ;
      RECT  4.545000  1.035000  4.785000 1.905000 ;
      RECT  4.685000  2.190000  5.755000 2.360000 ;
      RECT  4.725000  0.365000  5.465000 0.535000 ;
      RECT  4.975000  1.655000  5.415000 2.010000 ;
      RECT  5.295000  0.535000  5.465000 1.315000 ;
      RECT  5.295000  1.315000  6.095000 1.485000 ;
      RECT  5.585000  1.485000  6.095000 1.575000 ;
      RECT  5.585000  1.575000  5.755000 2.190000 ;
      RECT  5.635000  0.765000  6.435000 1.065000 ;
      RECT  5.635000  1.065000  5.805000 1.095000 ;
      RECT  5.715000  0.085000  6.085000 0.585000 ;
      RECT  5.925000  1.245000  6.095000 1.315000 ;
      RECT  5.925000  1.835000  6.095000 2.635000 ;
      RECT  6.265000  0.365000  6.725000 0.535000 ;
      RECT  6.265000  0.535000  6.435000 0.765000 ;
      RECT  6.265000  1.065000  6.435000 2.135000 ;
      RECT  6.265000  2.135000  6.515000 2.465000 ;
      RECT  6.605000  0.705000  7.155000 1.035000 ;
      RECT  6.605000  1.245000  6.795000 1.965000 ;
      RECT  6.740000  2.165000  7.625000 2.335000 ;
      RECT  6.955000  0.365000  7.495000 0.535000 ;
      RECT  6.965000  1.035000  7.155000 1.575000 ;
      RECT  6.965000  1.575000  7.285000 1.905000 ;
      RECT  7.325000  0.535000  7.495000 0.995000 ;
      RECT  7.325000  0.995000  8.370000 1.325000 ;
      RECT  7.325000  1.325000  7.625000 1.405000 ;
      RECT  7.455000  1.405000  7.625000 2.165000 ;
      RECT  7.740000  0.085000  8.110000 0.615000 ;
      RECT  7.795000  1.575000  8.725000 1.905000 ;
      RECT  7.805000  2.135000  8.110000 2.635000 ;
      RECT  8.360000  0.300000  8.725000 0.825000 ;
      RECT  8.395000  1.905000  8.725000 2.455000 ;
      RECT  8.540000  0.825000  8.725000 0.995000 ;
      RECT  8.540000  0.995000  9.275000 1.325000 ;
      RECT  8.540000  1.325000  8.725000 1.575000 ;
      RECT  8.895000  0.085000  9.085000 0.695000 ;
      RECT  8.895000  1.625000  9.075000 2.635000 ;
      RECT  9.755000  0.085000  9.985000 0.690000 ;
      RECT  9.765000  1.615000  9.935000 2.635000 ;
      RECT 10.205000  0.345000 10.455000 0.995000 ;
      RECT 10.205000  0.995000 11.065000 1.325000 ;
      RECT 10.205000  1.325000 10.535000 2.425000 ;
      RECT 10.690000  0.085000 11.020000 0.805000 ;
      RECT 10.715000  1.495000 11.020000 2.635000 ;
      RECT 11.610000  0.085000 11.780000 0.955000 ;
      RECT 11.610000  1.395000 11.780000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.645000  1.785000  0.815000 1.955000 ;
      RECT  1.050000  0.765000  1.220000 0.935000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  0.765000  4.915000 0.935000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.625000  1.785000  6.795000 1.955000 ;
      RECT  6.640000  0.765000  6.810000 0.935000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 6.855000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 0.990000 0.735000 1.280000 0.780000 ;
      RECT 0.990000 0.780000 6.870000 0.920000 ;
      RECT 0.990000 0.920000 1.280000 0.965000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 6.565000 1.755000 6.855000 1.800000 ;
      RECT 6.565000 1.940000 6.855000 1.985000 ;
      RECT 6.580000 0.735000 6.870000 0.780000 ;
      RECT 6.580000 0.920000 6.870000 0.965000 ;
  END
END sky130_fd_sc_hd__sdfxbp_2
MACRO sky130_fd_sc_hd__fahcin_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fahcin_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.42000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 1.075000 1.340000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.691500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 0.665000 1.740000 1.325000 ;
      LAYER mcon ;
        RECT 1.525000 0.765000 1.695000 0.935000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.240000 0.645000 4.490000 1.325000 ;
      LAYER mcon ;
        RECT 4.285000 0.765000 4.455000 0.935000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465000 0.735000 1.755000 0.780000 ;
        RECT 1.465000 0.780000 4.515000 0.920000 ;
        RECT 1.465000 0.920000 1.755000 0.965000 ;
        RECT 4.225000 0.735000 4.515000 0.780000 ;
        RECT 4.225000 0.920000 4.515000 0.965000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.493500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.520000 1.075000 10.965000 1.275000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.402800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.600000 0.755000 6.925000 0.925000 ;
        RECT 6.600000 0.925000 6.870000 1.675000 ;
        RECT 6.700000 1.675000 6.870000 1.785000 ;
        RECT 6.755000 0.595000 6.925000 0.755000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.470250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995000 0.255000 12.335000 0.825000 ;
        RECT 12.000000 1.785000 12.335000 2.465000 ;
        RECT 12.125000 0.825000 12.335000 1.785000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 12.420000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.610000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 12.420000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.420000 0.085000 ;
      RECT  0.000000  2.635000 12.420000 2.805000 ;
      RECT  0.085000  0.735000  0.430000 0.805000 ;
      RECT  0.085000  0.805000  0.255000 1.500000 ;
      RECT  0.085000  1.500000  0.440000 1.840000 ;
      RECT  0.085000  1.840000  1.110000 2.010000 ;
      RECT  0.085000  2.010000  0.430000 2.465000 ;
      RECT  0.100000  0.255000  0.430000 0.735000 ;
      RECT  0.425000  0.995000  0.780000 1.325000 ;
      RECT  0.600000  2.180000  0.770000 2.635000 ;
      RECT  0.610000  0.735000  1.325000 0.905000 ;
      RECT  0.610000  0.905000  0.780000 0.995000 ;
      RECT  0.610000  1.325000  0.780000 1.500000 ;
      RECT  0.610000  1.500000  1.450000 1.670000 ;
      RECT  0.630000  0.085000  0.800000 0.545000 ;
      RECT  0.940000  2.010000  1.110000 2.215000 ;
      RECT  0.940000  2.215000  1.970000 2.295000 ;
      RECT  0.940000  2.295000  3.515000 2.385000 ;
      RECT  0.995000  0.255000  3.390000 0.425000 ;
      RECT  0.995000  0.425000  2.100000 0.465000 ;
      RECT  0.995000  0.465000  1.325000 0.735000 ;
      RECT  1.280000  1.670000  1.450000 1.785000 ;
      RECT  1.280000  1.785000  2.050000 1.955000 ;
      RECT  1.280000  1.955000  1.450000 2.045000 ;
      RECT  1.715000  2.385000  3.515000 2.465000 ;
      RECT  1.985000  0.675000  2.390000 1.350000 ;
      RECT  2.220000  0.595000  2.390000 0.675000 ;
      RECT  2.220000  1.350000  2.390000 1.785000 ;
      RECT  2.515000  0.425000  3.390000 0.465000 ;
      RECT  2.565000  1.785000  2.895000 2.045000 ;
      RECT  2.620000  0.655000  3.025000 0.735000 ;
      RECT  2.620000  0.735000  3.135000 0.755000 ;
      RECT  2.620000  0.755000  3.730000 0.905000 ;
      RECT  2.640000  1.075000  2.970000 1.095000 ;
      RECT  2.640000  1.095000  3.120000 1.245000 ;
      RECT  2.800000  1.245000  3.120000 1.265000 ;
      RECT  2.950000  1.265000  3.120000 1.615000 ;
      RECT  3.055000  0.905000  3.730000 0.925000 ;
      RECT  3.215000  0.465000  3.390000 0.585000 ;
      RECT  3.245000  2.110000  3.460000 2.295000 ;
      RECT  3.290000  0.925000  3.460000 2.110000 ;
      RECT  3.560000  0.255000  4.570000 0.425000 ;
      RECT  3.560000  0.425000  3.730000 0.755000 ;
      RECT  3.710000  1.150000  4.070000 1.320000 ;
      RECT  3.710000  1.320000  3.880000 2.290000 ;
      RECT  3.710000  2.290000  5.065000 2.460000 ;
      RECT  3.900000  0.595000  4.070000 1.150000 ;
      RECT  4.080000  1.695000  4.445000 2.120000 ;
      RECT  4.240000  0.425000  4.570000 0.475000 ;
      RECT  4.690000  1.385000  5.170000 1.725000 ;
      RECT  4.815000  1.895000  5.995000 2.065000 ;
      RECT  4.815000  2.065000  5.065000 2.290000 ;
      RECT  4.830000  0.510000  5.000000 0.995000 ;
      RECT  4.830000  0.995000  5.630000 1.325000 ;
      RECT  4.830000  1.325000  5.170000 1.385000 ;
      RECT  5.180000  0.085000  5.510000 0.805000 ;
      RECT  5.260000  2.235000  5.590000 2.635000 ;
      RECT  5.635000  1.555000  6.370000 1.725000 ;
      RECT  5.680000  0.380000  5.970000 0.815000 ;
      RECT  5.800000  0.815000  5.970000 1.555000 ;
      RECT  5.825000  2.065000  5.995000 2.295000 ;
      RECT  5.825000  2.295000  7.950000 2.465000 ;
      RECT  6.140000  0.740000  6.425000 1.325000 ;
      RECT  6.200000  1.725000  6.370000 1.895000 ;
      RECT  6.200000  1.895000  6.530000 1.955000 ;
      RECT  6.200000  1.955000  7.210000 2.125000 ;
      RECT  6.255000  0.255000  7.695000 0.425000 ;
      RECT  6.255000  0.425000  6.585000 0.570000 ;
      RECT  7.040000  1.060000  7.270000 1.230000 ;
      RECT  7.040000  1.230000  7.210000 1.955000 ;
      RECT  7.100000  0.595000  7.350000 0.925000 ;
      RECT  7.100000  0.925000  7.270000 1.060000 ;
      RECT  7.380000  1.360000  7.610000 1.530000 ;
      RECT  7.380000  1.530000  7.550000 2.125000 ;
      RECT  7.440000  1.105000  7.695000 1.290000 ;
      RECT  7.440000  1.290000  7.610000 1.360000 ;
      RECT  7.520000  0.425000  7.695000 1.105000 ;
      RECT  7.780000  1.550000  8.035000 1.720000 ;
      RECT  7.780000  1.720000  7.950000 2.295000 ;
      RECT  7.865000  0.255000  9.980000 0.425000 ;
      RECT  7.865000  0.425000  8.035000 0.740000 ;
      RECT  7.865000  0.995000  8.035000 1.550000 ;
      RECT  8.220000  1.955000  8.390000 2.295000 ;
      RECT  8.220000  2.295000  9.410000 2.465000 ;
      RECT  8.305000  0.595000  8.555000 0.925000 ;
      RECT  8.375000  0.925000  8.555000 1.445000 ;
      RECT  8.375000  1.445000  8.670000 1.530000 ;
      RECT  8.375000  1.530000  8.890000 1.785000 ;
      RECT  8.560000  1.785000  8.890000 2.125000 ;
      RECT  8.725000  0.595000  9.410000 0.765000 ;
      RECT  8.835000  0.995000  9.070000 1.325000 ;
      RECT  9.240000  0.765000  9.410000 1.875000 ;
      RECT  9.240000  1.875000 10.885000 2.025000 ;
      RECT  9.240000  2.025000 10.145000 2.030000 ;
      RECT  9.240000  2.030000 10.130000 2.035000 ;
      RECT  9.240000  2.035000 10.120000 2.040000 ;
      RECT  9.240000  2.040000 10.105000 2.045000 ;
      RECT  9.240000  2.045000  9.410000 2.295000 ;
      RECT  9.640000  0.425000  9.980000 0.825000 ;
      RECT  9.640000  0.825000  9.810000 1.535000 ;
      RECT  9.640000  1.535000 10.010000 1.705000 ;
      RECT  9.980000  0.995000 10.350000 1.325000 ;
      RECT 10.055000  1.870000 10.885000 1.875000 ;
      RECT 10.070000  1.865000 10.885000 1.870000 ;
      RECT 10.085000  1.860000 10.885000 1.865000 ;
      RECT 10.100000  1.855000 10.885000 1.860000 ;
      RECT 10.180000  0.085000 10.350000 0.565000 ;
      RECT 10.180000  0.735000 10.910000 0.905000 ;
      RECT 10.180000  0.905000 10.350000 0.995000 ;
      RECT 10.180000  1.325000 10.350000 1.445000 ;
      RECT 10.180000  1.445000 10.885000 1.855000 ;
      RECT 10.190000  2.195000 10.360000 2.635000 ;
      RECT 10.530000  0.285000 10.910000 0.735000 ;
      RECT 10.535000  2.025000 10.885000 2.465000 ;
      RECT 11.075000  1.455000 11.405000 2.465000 ;
      RECT 11.155000  0.270000 11.325000 0.680000 ;
      RECT 11.155000  0.680000 11.405000 1.455000 ;
      RECT 11.495000  0.085000 11.825000 0.510000 ;
      RECT 11.575000  1.785000 11.830000 2.635000 ;
      RECT 11.645000  0.995000 11.955000 1.615000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.880000  1.785000  2.050000 1.955000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  1.105000  2.155000 1.275000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.570000  1.785000  2.740000 1.955000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  2.950000  1.445000  3.120000 1.615000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.140000  1.785000  4.310000 1.955000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.760000  1.445000  4.930000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.140000  1.105000  6.310000 1.275000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.520000  0.765000  7.690000 0.935000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.440000  1.445000  8.610000 1.615000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  8.900000  1.105000  9.070000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.220000  0.765000 11.390000 0.935000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 11.680000  1.445000 11.850000 1.615000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
    LAYER met1 ;
      RECT  1.820000 1.755000  2.110000 1.800000 ;
      RECT  1.820000 1.800000  4.370000 1.940000 ;
      RECT  1.820000 1.940000  2.110000 1.985000 ;
      RECT  1.925000 1.075000  2.215000 1.120000 ;
      RECT  1.925000 1.120000  9.130000 1.260000 ;
      RECT  1.925000 1.260000  2.215000 1.305000 ;
      RECT  2.510000 1.755000  2.800000 1.800000 ;
      RECT  2.510000 1.940000  2.800000 1.985000 ;
      RECT  2.890000 1.415000  3.180000 1.460000 ;
      RECT  2.890000 1.460000  4.990000 1.600000 ;
      RECT  2.890000 1.600000  3.180000 1.645000 ;
      RECT  4.080000 1.755000  4.370000 1.800000 ;
      RECT  4.080000 1.940000  4.370000 1.985000 ;
      RECT  4.700000 1.415000  4.990000 1.460000 ;
      RECT  4.700000 1.600000  4.990000 1.645000 ;
      RECT  6.080000 1.075000  6.370000 1.120000 ;
      RECT  6.080000 1.260000  6.370000 1.305000 ;
      RECT  7.460000 0.735000  7.750000 0.780000 ;
      RECT  7.460000 0.780000 11.450000 0.920000 ;
      RECT  7.460000 0.920000  7.750000 0.965000 ;
      RECT  8.380000 1.415000  8.670000 1.460000 ;
      RECT  8.380000 1.460000 11.910000 1.600000 ;
      RECT  8.380000 1.600000  8.670000 1.645000 ;
      RECT  8.840000 1.075000  9.130000 1.120000 ;
      RECT  8.840000 1.260000  9.130000 1.305000 ;
      RECT 11.160000 0.735000 11.450000 0.780000 ;
      RECT 11.160000 0.920000 11.450000 0.965000 ;
      RECT 11.620000 1.415000 11.910000 1.460000 ;
      RECT 11.620000 1.600000 11.910000 1.645000 ;
  END
END sky130_fd_sc_hd__fahcin_1
MACRO sky130_fd_sc_hd__sdfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfsbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.34000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.915000 0.275000 13.255000 0.825000 ;
        RECT 12.915000 1.495000 13.255000 2.450000 ;
        RECT 13.070000 0.825000 13.255000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.500000 0.255000 11.830000 2.465000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.345000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.765000 0.825000 1.675000 ;
      LAYER mcon ;
        RECT 0.610000 1.105000 0.780000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.370000 1.075000 2.700000 1.600000 ;
      LAYER mcon ;
        RECT 2.445000 1.105000 2.615000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.550000 1.075000 0.840000 1.120000 ;
        RECT 0.550000 1.120000 2.675000 1.260000 ;
        RECT 0.550000 1.260000 0.840000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.015000 1.765000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.885000 1.415000  9.110000 1.525000 ;
        RECT 8.885000 1.525000 10.075000 1.725000 ;
      LAYER mcon ;
        RECT 8.885000 1.445000 9.055000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.115000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.825000 1.415000 9.115000 1.460000 ;
        RECT 8.825000 1.600000 9.115000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.590000 ;
        RECT 2.905000 1.590000 3.085000 1.960000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 13.530000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.340000 0.085000 ;
      RECT  0.000000  2.635000 13.340000 2.805000 ;
      RECT  0.085000  0.085000  0.480000 0.595000 ;
      RECT  0.085000  1.845000  1.105000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.765000 2.635000 ;
      RECT  0.875000  0.280000  1.655000 0.560000 ;
      RECT  0.935000  2.025000  1.105000 2.255000 ;
      RECT  0.935000  2.255000  2.045000 2.465000 ;
      RECT  1.295000  1.870000  1.695000 2.075000 ;
      RECT  1.380000  0.560000  1.655000 0.590000 ;
      RECT  1.380000  0.590000  1.660000 0.600000 ;
      RECT  1.395000  0.600000  1.660000 0.605000 ;
      RECT  1.405000  0.605000  1.660000 0.610000 ;
      RECT  1.420000  0.610000  1.660000 0.615000 ;
      RECT  1.430000  0.615000  1.670000 0.620000 ;
      RECT  1.440000  0.620000  1.670000 0.630000 ;
      RECT  1.445000  0.630000  1.670000 0.635000 ;
      RECT  1.460000  0.635000  1.670000 0.645000 ;
      RECT  1.475000  0.645000  1.670000 0.655000 ;
      RECT  1.475000  0.655000  1.695000 0.665000 ;
      RECT  1.495000  0.665000  1.695000 0.705000 ;
      RECT  1.505000  0.705000  1.695000 1.870000 ;
      RECT  1.825000  0.085000  2.005000 0.545000 ;
      RECT  1.865000  0.715000  2.515000 0.905000 ;
      RECT  1.865000  0.905000  2.200000 1.770000 ;
      RECT  1.865000  1.770000  2.520000 2.085000 ;
      RECT  2.260000  0.255000  2.515000 0.715000 ;
      RECT  2.270000  2.085000  2.520000 2.465000 ;
      RECT  2.690000  0.085000  3.030000 0.555000 ;
      RECT  2.690000  2.140000  3.030000 2.635000 ;
      RECT  3.255000  1.775000  3.995000 1.955000 ;
      RECT  3.255000  1.955000  3.425000 2.325000 ;
      RECT  3.270000  0.255000  3.455000 0.715000 ;
      RECT  3.270000  0.715000  3.995000 0.885000 ;
      RECT  3.595000  2.275000  3.925000 2.635000 ;
      RECT  3.630000  0.085000  3.940000 0.545000 ;
      RECT  3.735000  0.885000  3.995000 1.775000 ;
      RECT  4.095000  2.135000  4.440000 2.465000 ;
      RECT  4.110000  0.255000  4.335000 0.585000 ;
      RECT  4.165000  0.585000  4.335000 1.090000 ;
      RECT  4.165000  1.090000  4.490000 1.420000 ;
      RECT  4.165000  1.420000  4.440000 2.135000 ;
      RECT  4.505000  0.255000  4.830000 0.920000 ;
      RECT  4.610000  1.590000  4.915000 1.615000 ;
      RECT  4.610000  1.615000  4.830000 2.465000 ;
      RECT  4.660000  0.920000  4.830000 1.445000 ;
      RECT  4.660000  1.445000  4.915000 1.590000 ;
      RECT  5.000000  0.255000  5.440000 1.225000 ;
      RECT  5.000000  1.225000  7.660000 1.275000 ;
      RECT  5.030000  2.135000  5.755000 2.465000 ;
      RECT  5.085000  1.275000  6.435000 1.395000 ;
      RECT  5.205000  1.575000  5.415000 1.955000 ;
      RECT  5.585000  1.395000  5.755000 2.135000 ;
      RECT  5.610000  0.085000  6.095000 0.465000 ;
      RECT  5.610000  0.635000  6.535000 0.805000 ;
      RECT  5.610000  0.805000  5.975000 1.015000 ;
      RECT  5.925000  1.575000  6.095000 1.935000 ;
      RECT  5.925000  1.935000  6.765000 2.105000 ;
      RECT  5.945000  2.275000  6.275000 2.635000 ;
      RECT  6.250000  0.975000  7.660000 1.225000 ;
      RECT  6.275000  0.255000  6.535000 0.635000 ;
      RECT  6.550000  2.105000  6.765000 2.450000 ;
      RECT  6.735000  0.085000  7.630000 0.805000 ;
      RECT  7.005000  2.125000  7.960000 2.635000 ;
      RECT  7.190000  1.495000  8.005000 1.955000 ;
      RECT  7.300000  1.275000  7.660000 1.325000 ;
      RECT  7.835000  0.695000  9.040000 0.895000 ;
      RECT  7.835000  0.895000  8.005000 1.495000 ;
      RECT  8.130000  2.125000  8.935000 2.460000 ;
      RECT  8.365000  1.075000  8.595000 1.905000 ;
      RECT  8.410000  0.275000  9.825000 0.445000 ;
      RECT  8.765000  1.895000 10.465000 2.065000 ;
      RECT  8.765000  2.065000  8.935000 2.125000 ;
      RECT  8.810000  0.895000  9.040000 1.245000 ;
      RECT  9.195000  2.235000  9.525000 2.635000 ;
      RECT  9.290000  0.855000  9.465000 1.185000 ;
      RECT  9.290000  1.185000 10.895000 1.355000 ;
      RECT  9.655000  0.445000  9.825000 0.845000 ;
      RECT  9.655000  0.845000 10.545000 1.015000 ;
      RECT  9.695000  2.065000  9.910000 2.450000 ;
      RECT 10.135000  2.235000 10.465000 2.635000 ;
      RECT 10.220000  0.085000 10.390000 0.545000 ;
      RECT 10.245000  1.525000 10.465000 1.895000 ;
      RECT 10.560000  0.255000 10.895000 0.540000 ;
      RECT 10.635000  1.355000 10.895000 2.465000 ;
      RECT 10.715000  0.540000 10.895000 1.185000 ;
      RECT 11.120000  0.085000 11.330000 0.885000 ;
      RECT 11.120000  1.485000 11.330000 2.635000 ;
      RECT 12.060000  0.255000 12.270000 0.995000 ;
      RECT 12.060000  0.995000 12.900000 1.325000 ;
      RECT 12.060000  1.325000 12.270000 2.465000 ;
      RECT 12.540000  0.085000 12.745000 0.825000 ;
      RECT 12.575000  1.575000 12.745000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.445000  1.695000 1.615000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  1.785000  3.995000 1.955000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.445000  4.915000 1.615000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  1.785000  5.375000 1.955000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  1.785000  7.675000 1.955000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  1.105000  8.595000 1.275000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.975000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.735000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.655000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.685000 1.415000 4.975000 1.460000 ;
      RECT 4.685000 1.600000 4.975000 1.645000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 7.445000 1.755000 7.735000 1.800000 ;
      RECT 7.445000 1.940000 7.735000 1.985000 ;
      RECT 8.365000 1.075000 8.655000 1.120000 ;
      RECT 8.365000 1.260000 8.655000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfsbp_1
MACRO sky130_fd_sc_hd__sdfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfsbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.26000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.410000 0.275000 13.740000 0.825000 ;
        RECT 13.410000 1.495000 13.740000 2.450000 ;
        RECT 13.515000 0.825000 13.740000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.460000 0.255000 11.855000 2.465000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.765000 0.820000 1.675000 ;
      LAYER mcon ;
        RECT 0.605000 1.105000 0.775000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.405000 1.075000 2.735000 1.590000 ;
      LAYER mcon ;
        RECT 2.445000 1.105000 2.615000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545000 1.075000 0.835000 1.120000 ;
        RECT 0.545000 1.120000 2.675000 1.260000 ;
        RECT 0.545000 1.260000 0.835000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.065000 1.765000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.880000 1.435000 9.115000 1.525000 ;
        RECT 8.880000 1.525000 9.935000 1.725000 ;
      LAYER mcon ;
        RECT 8.940000 1.445000 9.110000 1.615000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.170000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.880000 1.415000 9.170000 1.460000 ;
        RECT 8.880000 1.600000 9.170000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.615000 ;
        RECT 2.905000 1.615000 3.100000 1.970000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 14.450000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.260000 0.085000 ;
      RECT  0.000000  2.635000 14.260000 2.805000 ;
      RECT  0.085000  0.085000  0.700000 0.595000 ;
      RECT  0.085000  1.845000  1.185000 2.075000 ;
      RECT  0.085000  2.075000  0.345000 2.465000 ;
      RECT  0.515000  2.275000  0.845000 2.635000 ;
      RECT  0.870000  0.255000  1.670000 0.595000 ;
      RECT  1.015000  2.075000  1.185000 2.255000 ;
      RECT  1.015000  2.255000  2.105000 2.465000 ;
      RECT  1.355000  1.845000  1.695000 2.085000 ;
      RECT  1.495000  0.595000  1.670000 0.645000 ;
      RECT  1.495000  0.645000  1.695000 0.705000 ;
      RECT  1.500000  0.705000  1.695000 0.720000 ;
      RECT  1.505000  0.720000  1.695000 1.845000 ;
      RECT  1.840000  0.085000  2.090000 0.545000 ;
      RECT  1.980000  0.715000  2.530000 0.905000 ;
      RECT  1.980000  0.905000  2.235000 1.760000 ;
      RECT  1.980000  1.760000  2.535000 2.085000 ;
      RECT  2.260000  0.255000  2.530000 0.715000 ;
      RECT  2.275000  2.085000  2.535000 2.465000 ;
      RECT  2.700000  0.085000  3.100000 0.555000 ;
      RECT  2.705000  2.140000  3.100000 2.635000 ;
      RECT  3.270000  0.255000  3.470000 0.715000 ;
      RECT  3.270000  0.715000  3.995000 0.885000 ;
      RECT  3.270000  1.830000  3.995000 2.000000 ;
      RECT  3.270000  2.000000  3.475000 2.325000 ;
      RECT  3.640000  0.085000  3.940000 0.545000 ;
      RECT  3.645000  2.275000  3.975000 2.635000 ;
      RECT  3.735000  0.885000  3.995000 1.830000 ;
      RECT  4.110000  0.255000  4.335000 0.585000 ;
      RECT  4.145000  2.135000  4.440000 2.465000 ;
      RECT  4.165000  0.585000  4.335000 1.090000 ;
      RECT  4.165000  1.090000  4.490000 1.420000 ;
      RECT  4.165000  1.420000  4.440000 2.135000 ;
      RECT  4.505000  0.255000  4.885000 0.920000 ;
      RECT  4.665000  1.590000  4.970000 1.615000 ;
      RECT  4.665000  1.615000  4.890000 2.465000 ;
      RECT  4.715000  0.920000  4.885000 1.445000 ;
      RECT  4.715000  1.445000  4.970000 1.590000 ;
      RECT  5.055000  0.255000  5.450000 1.225000 ;
      RECT  5.055000  1.225000  7.705000 1.275000 ;
      RECT  5.060000  2.135000  5.805000 2.465000 ;
      RECT  5.140000  1.275000  6.475000 1.395000 ;
      RECT  5.205000  1.575000  5.465000 1.955000 ;
      RECT  5.620000  0.635000  6.550000 0.805000 ;
      RECT  5.620000  0.805000  6.015000 1.015000 ;
      RECT  5.635000  1.395000  5.805000 2.135000 ;
      RECT  5.665000  0.085000  6.165000 0.465000 ;
      RECT  5.975000  1.575000  6.145000 1.935000 ;
      RECT  5.975000  1.935000  6.820000 2.105000 ;
      RECT  6.000000  2.275000  6.330000 2.635000 ;
      RECT  6.305000  0.975000  7.705000 1.225000 ;
      RECT  6.335000  0.255000  6.550000 0.635000 ;
      RECT  6.605000  2.105000  6.820000 2.450000 ;
      RECT  6.720000  0.085000  7.705000 0.805000 ;
      RECT  7.060000  2.125000  8.015000 2.635000 ;
      RECT  7.355000  1.275000  7.705000 1.325000 ;
      RECT  7.385000  1.705000  8.055000 1.955000 ;
      RECT  7.885000  0.695000  9.085000 0.895000 ;
      RECT  7.885000  0.895000  8.055000 1.705000 ;
      RECT  8.185000  2.125000  8.990000 2.460000 ;
      RECT  8.420000  1.075000  8.650000 1.905000 ;
      RECT  8.465000  0.275000  9.855000 0.515000 ;
      RECT  8.820000  1.895000 10.430000 2.065000 ;
      RECT  8.820000  2.065000  8.990000 2.125000 ;
      RECT  8.830000  0.895000  9.085000 1.265000 ;
      RECT  9.160000  2.235000  9.490000 2.635000 ;
      RECT  9.285000  0.855000  9.515000 1.185000 ;
      RECT  9.285000  1.185000 10.910000 1.355000 ;
      RECT  9.660000  2.065000  9.930000 2.450000 ;
      RECT  9.685000  0.515000  9.855000 0.845000 ;
      RECT  9.685000  0.845000 10.560000 1.015000 ;
      RECT 10.035000  0.085000 10.285000 0.545000 ;
      RECT 10.100000  2.235000 10.430000 2.635000 ;
      RECT 10.105000  1.525000 10.430000 1.895000 ;
      RECT 10.465000  0.255000 10.910000 0.585000 ;
      RECT 10.600000  1.355000 10.845000 2.465000 ;
      RECT 10.730000  0.585000 10.910000 1.185000 ;
      RECT 11.080000  1.485000 11.290000 2.635000 ;
      RECT 11.120000  0.085000 11.290000 0.885000 ;
      RECT 12.025000  0.085000 12.315000 0.885000 ;
      RECT 12.025000  1.485000 12.315000 2.635000 ;
      RECT 12.530000  0.255000 12.715000 0.995000 ;
      RECT 12.530000  0.995000 13.345000 1.325000 ;
      RECT 12.530000  1.325000 12.715000 2.465000 ;
      RECT 12.885000  0.085000 13.240000 0.825000 ;
      RECT 12.885000  1.635000 13.240000 2.635000 ;
      RECT 13.910000  0.085000 14.175000 0.885000 ;
      RECT 13.910000  1.485000 14.175000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.445000  1.695000 1.615000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  1.785000  3.995000 1.955000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  1.105000  4.455000 1.275000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  4.800000  1.445000  4.970000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.260000  1.785000  5.430000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.560000  1.785000  7.730000 1.955000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.480000  1.105000  8.650000 1.275000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 5.030000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.790000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.710000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.740000 1.415000 5.030000 1.460000 ;
      RECT 4.740000 1.600000 5.030000 1.645000 ;
      RECT 5.200000 1.755000 5.490000 1.800000 ;
      RECT 5.200000 1.940000 5.490000 1.985000 ;
      RECT 7.500000 1.755000 7.790000 1.800000 ;
      RECT 7.500000 1.940000 7.790000 1.985000 ;
      RECT 8.420000 1.075000 8.710000 1.120000 ;
      RECT 8.420000 1.260000 8.710000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfsbp_2
MACRO sky130_fd_sc_hd__nor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.810000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.980000 1.075000 1.750000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 1.705000 0.735000 ;
        RECT 0.535000 0.735000 2.135000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 1.375000 1.445000 2.135000 1.665000 ;
        RECT 1.375000 1.665000 1.705000 2.125000 ;
        RECT 1.920000 0.905000 2.135000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 1.205000 1.665000 ;
      RECT 0.090000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.865000 2.635000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.035000  1.665000 1.205000 2.295000 ;
      RECT 1.035000  2.295000 2.175000 2.465000 ;
      RECT 1.875000  0.085000 2.165000 0.555000 ;
      RECT 1.875000  1.835000 2.175000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2_2
MACRO sky130_fd_sc_hd__nor2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.360000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.075000 3.530000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.800000 1.075000 6.540000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 7.275000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 3.895000 0.255000 4.225000 0.725000 ;
        RECT 3.935000 1.445000 7.275000 1.615000 ;
        RECT 3.935000 1.615000 4.185000 2.125000 ;
        RECT 4.735000 0.255000 5.065000 0.725000 ;
        RECT 4.775000 1.615000 5.025000 2.125000 ;
        RECT 5.575000 0.255000 5.905000 0.725000 ;
        RECT 5.615000 1.615000 5.865000 2.125000 ;
        RECT 6.415000 0.255000 6.745000 0.725000 ;
        RECT 6.455000 1.615000 6.705000 2.125000 ;
        RECT 6.710000 0.905000 7.275000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 7.550000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 3.765000 1.665000 ;
      RECT 0.090000  1.665000 0.405000 2.465000 ;
      RECT 0.575000  1.835000 0.825000 2.635000 ;
      RECT 0.995000  1.665000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.835000 1.665000 2.635000 ;
      RECT 1.835000  1.665000 2.085000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.255000  1.835000 2.505000 2.635000 ;
      RECT 2.675000  1.665000 2.925000 2.465000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 3.095000  1.835000 3.345000 2.635000 ;
      RECT 3.515000  1.665000 3.765000 2.295000 ;
      RECT 3.515000  2.295000 7.125000 2.465000 ;
      RECT 3.555000  0.085000 3.725000 0.555000 ;
      RECT 4.355000  1.785000 4.605000 2.295000 ;
      RECT 4.395000  0.085000 4.565000 0.555000 ;
      RECT 5.195000  1.785000 5.445000 2.295000 ;
      RECT 5.235000  0.085000 5.405000 0.555000 ;
      RECT 6.035000  1.785000 6.285000 2.295000 ;
      RECT 6.075000  0.085000 6.245000 0.555000 ;
      RECT 6.875000  1.785000 7.125000 2.295000 ;
      RECT 6.915000  0.085000 7.205000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2_8
MACRO sky130_fd_sc_hd__nor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 1.075000 1.295000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.435000 1.325000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.495000 0.775000 1.665000 ;
        RECT 0.095000 1.665000 0.425000 2.450000 ;
        RECT 0.515000 0.255000 0.845000 0.895000 ;
        RECT 0.605000 0.895000 0.775000 1.495000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 1.570000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.380000 0.085000 ;
      RECT 0.000000  2.635000 1.380000 2.805000 ;
      RECT 0.105000  0.085000 0.345000 0.895000 ;
      RECT 0.955000  1.495000 1.285000 2.635000 ;
      RECT 1.015000  0.085000 1.285000 0.895000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2_1
MACRO sky130_fd_sc_hd__nor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.800000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.120000 1.075000 3.485000 1.275000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 4.055000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 2.295000 1.445000 4.055000 1.745000 ;
        RECT 2.295000 1.745000 2.465000 2.125000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 3.135000 1.745000 3.305000 2.125000 ;
        RECT 3.655000 0.905000 4.055000 1.445000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 2.125000 1.665000 ;
      RECT 0.090000  1.665000 0.365000 2.465000 ;
      RECT 0.535000  1.835000 0.865000 2.635000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.035000  1.665000 1.205000 2.465000 ;
      RECT 1.375000  1.835000 1.625000 2.635000 ;
      RECT 1.795000  1.665000 2.125000 2.295000 ;
      RECT 1.795000  2.295000 3.890000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.635000  1.935000 2.965000 2.295000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 3.475000  1.915000 3.890000 2.295000 ;
      RECT 3.555000  0.085000 3.840000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
END sky130_fd_sc_hd__nor2_4
MACRO sky130_fd_sc_hd__nor4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.180000 1.075000 1.825000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095000 1.075000 4.070000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.295000 1.075000 5.705000 1.285000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.875000 1.075000 7.295000 1.285000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 7.735000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.215000 0.255000 2.545000 0.725000 ;
        RECT 3.055000 0.255000 3.385000 0.725000 ;
        RECT 4.415000 0.255000 4.745000 0.725000 ;
        RECT 5.255000 0.255000 5.585000 0.725000 ;
        RECT 6.095000 0.255000 6.425000 0.725000 ;
        RECT 6.135000 1.455000 7.735000 1.625000 ;
        RECT 6.135000 1.625000 6.385000 2.125000 ;
        RECT 6.935000 0.255000 7.265000 0.725000 ;
        RECT 6.975000 1.625000 7.225000 2.125000 ;
        RECT 7.465000 0.905000 7.735000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 2.085000 1.625000 ;
      RECT 0.090000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.995000  1.625000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.795000 1.665000 2.635000 ;
      RECT 1.835000  1.625000 2.085000 2.295000 ;
      RECT 1.835000  2.295000 3.820000 2.465000 ;
      RECT 1.875000  0.085000 2.045000 0.555000 ;
      RECT 2.255000  1.455000 5.545000 1.625000 ;
      RECT 2.255000  1.625000 2.505000 2.125000 ;
      RECT 2.675000  1.795000 2.925000 2.295000 ;
      RECT 2.715000  0.085000 2.885000 0.555000 ;
      RECT 3.095000  1.625000 3.345000 2.125000 ;
      RECT 3.515000  1.795000 3.820000 2.295000 ;
      RECT 3.555000  0.085000 4.245000 0.555000 ;
      RECT 4.005000  1.795000 4.285000 2.295000 ;
      RECT 4.005000  2.295000 7.645000 2.465000 ;
      RECT 4.455000  1.625000 4.705000 2.125000 ;
      RECT 4.875000  1.795000 5.125000 2.295000 ;
      RECT 4.915000  0.085000 5.085000 0.555000 ;
      RECT 5.295000  1.625000 5.545000 2.125000 ;
      RECT 5.715000  1.795000 5.965000 2.295000 ;
      RECT 5.755000  0.085000 5.925000 0.555000 ;
      RECT 6.555000  1.795000 6.805000 2.295000 ;
      RECT 6.595000  0.085000 6.765000 0.555000 ;
      RECT 7.395000  1.795000 7.645000 2.295000 ;
      RECT 7.435000  0.085000 7.605000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4_4
MACRO sky130_fd_sc_hd__nor4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.300000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 0.655000 2.215000 1.665000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245000 1.075000 1.695000 1.245000 ;
        RECT 1.455000 1.245000 1.695000 2.450000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845000 0.995000 1.075000 1.415000 ;
        RECT 0.845000 1.415000 1.285000 1.615000 ;
        RECT 1.030000 1.615000 1.285000 2.450000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.745000 0.335000 1.325000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.672750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.495000 0.675000 1.665000 ;
        RECT 0.090000 1.665000 0.425000 2.450000 ;
        RECT 0.505000 0.645000 0.860000 0.655000 ;
        RECT 0.505000 0.655000 1.705000 0.825000 ;
        RECT 0.505000 0.825000 0.675000 1.495000 ;
        RECT 0.595000 0.385000 0.860000 0.645000 ;
        RECT 1.535000 0.385000 1.705000 0.655000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.300000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 2.490000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.300000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.300000 0.085000 ;
      RECT 0.000000  2.635000 2.300000 2.805000 ;
      RECT 0.085000  0.085000 0.345000 0.575000 ;
      RECT 1.035000  0.085000 1.365000 0.485000 ;
      RECT 1.875000  0.085000 2.205000 0.485000 ;
      RECT 1.955000  1.835000 2.215000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4_1
MACRO sky130_fd_sc_hd__nor4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.200000 1.075000 0.965000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135000 1.075000 1.940000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.075000 3.105000 1.285000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.340000 1.075000 3.925000 1.285000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 4.515000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.775000 0.255000 3.105000 0.725000 ;
        RECT 3.615000 0.255000 3.945000 0.725000 ;
        RECT 3.655000 1.455000 4.515000 1.625000 ;
        RECT 3.655000 1.625000 3.905000 2.125000 ;
        RECT 4.180000 0.905000 4.515000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.150000  1.455000 2.085000 1.625000 ;
      RECT 0.150000  1.625000 0.405000 2.465000 ;
      RECT 0.575000  1.795000 0.825000 2.635000 ;
      RECT 0.995000  1.625000 1.245000 2.465000 ;
      RECT 1.035000  0.085000 1.205000 0.555000 ;
      RECT 1.415000  1.795000 1.665000 2.295000 ;
      RECT 1.415000  2.295000 3.065000 2.465000 ;
      RECT 1.835000  1.625000 2.085000 2.125000 ;
      RECT 1.875000  0.085000 2.605000 0.555000 ;
      RECT 2.395000  1.455000 3.485000 1.625000 ;
      RECT 2.395000  1.625000 2.645000 2.125000 ;
      RECT 2.815000  1.795000 3.065000 2.295000 ;
      RECT 3.235000  1.625000 3.485000 2.295000 ;
      RECT 3.235000  2.295000 4.325000 2.465000 ;
      RECT 3.275000  0.085000 3.445000 0.555000 ;
      RECT 4.075000  1.795000 4.325000 2.295000 ;
      RECT 4.115000  0.085000 4.405000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
END sky130_fd_sc_hd__nor4_2
MACRO sky130_fd_sc_hd__dlrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.060000 0.255000 6.410000 2.465000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.475000 0.255000 7.735000 0.595000 ;
        RECT 7.475000 1.785000 7.735000 2.465000 ;
        RECT 7.565000 0.595000 7.735000 1.785000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.450000 0.995000 5.435000 1.325000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.325000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.780000 0.805000 ;
      RECT 0.085000  1.795000 0.780000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 1.685000 ;
      RECT 2.600000  0.765000 3.095000 1.035000 ;
      RECT 2.745000  2.255000 3.585000 2.425000 ;
      RECT 2.770000  0.365000 3.500000 0.535000 ;
      RECT 2.925000  1.035000 3.095000 1.575000 ;
      RECT 2.925000  1.575000 3.265000 1.905000 ;
      RECT 2.925000  1.905000 3.130000 1.995000 ;
      RECT 3.270000  2.125000 3.585000 2.255000 ;
      RECT 3.305000  2.075000 3.585000 2.125000 ;
      RECT 3.330000  0.535000 3.500000 0.995000 ;
      RECT 3.330000  0.995000 4.200000 1.165000 ;
      RECT 3.395000  2.015000 3.605000 2.045000 ;
      RECT 3.395000  2.045000 3.585000 2.075000 ;
      RECT 3.415000  1.990000 3.605000 2.015000 ;
      RECT 3.420000  1.975000 3.605000 1.990000 ;
      RECT 3.430000  1.960000 3.605000 1.975000 ;
      RECT 3.435000  1.165000 4.200000 1.325000 ;
      RECT 3.435000  1.325000 3.605000 1.960000 ;
      RECT 3.735000  0.085000 4.070000 0.530000 ;
      RECT 3.755000  2.135000 4.590000 2.635000 ;
      RECT 3.840000  1.535000 5.890000 1.765000 ;
      RECT 3.840000  1.765000 4.950000 1.865000 ;
      RECT 4.240000  0.255000 4.540000 0.655000 ;
      RECT 4.240000  0.655000 5.890000 0.825000 ;
      RECT 4.780000  1.865000 4.950000 2.435000 ;
      RECT 5.120000  0.085000 5.890000 0.485000 ;
      RECT 5.120000  1.935000 5.890000 2.635000 ;
      RECT 5.655000  0.825000 5.890000 1.535000 ;
      RECT 6.580000  0.255000 6.805000 0.995000 ;
      RECT 6.580000  0.995000 7.395000 1.325000 ;
      RECT 6.580000  1.325000 6.830000 2.465000 ;
      RECT 6.975000  0.085000 7.305000 0.465000 ;
      RECT 7.010000  1.835000 7.305000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.445000 2.640000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.925000  1.785000 3.095000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 2.700000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 3.155000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.415000 2.700000 1.460000 ;
      RECT 2.410000 1.600000 2.700000 1.645000 ;
      RECT 2.865000 1.755000 3.155000 1.800000 ;
      RECT 2.865000 1.940000 3.155000 1.985000 ;
  END
END sky130_fd_sc_hd__dlrbp_1
MACRO sky130_fd_sc_hd__dlrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.460000 0.955000 1.790000 1.325000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.478500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.680000 0.330000 5.850000 0.665000 ;
        RECT 5.680000 0.665000 6.150000 0.835000 ;
        RECT 5.680000 1.495000 6.065000 1.660000 ;
        RECT 5.680000 1.660000 5.930000 2.465000 ;
        RECT 5.790000 0.835000 6.150000 0.885000 ;
        RECT 5.790000 0.885000 6.360000 1.325000 ;
        RECT 5.790000 1.325000 6.065000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.515000 0.255000 7.765000 0.825000 ;
        RECT 7.515000 1.605000 7.765000 2.465000 ;
        RECT 7.595000 0.825000 7.765000 1.055000 ;
        RECT 7.595000 1.055000 8.195000 1.325000 ;
        RECT 7.595000 1.325000 7.765000 1.605000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.400000 0.995000 5.150000 1.325000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.470000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.085000  0.345000 0.345000 0.635000 ;
      RECT 0.085000  0.635000 0.780000 0.805000 ;
      RECT 0.085000  1.795000 0.780000 1.965000 ;
      RECT 0.085000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.845000 0.465000 ;
      RECT 0.515000  2.135000 0.845000 2.635000 ;
      RECT 0.610000  0.805000 0.780000 1.070000 ;
      RECT 0.610000  1.070000 0.840000 1.400000 ;
      RECT 0.610000  1.400000 0.780000 1.795000 ;
      RECT 1.015000  0.345000 1.185000 1.685000 ;
      RECT 1.015000  1.685000 1.240000 2.465000 ;
      RECT 1.455000  1.495000 2.140000 1.665000 ;
      RECT 1.455000  1.665000 1.785000 2.415000 ;
      RECT 1.535000  0.345000 1.705000 0.615000 ;
      RECT 1.535000  0.615000 2.140000 0.765000 ;
      RECT 1.535000  0.765000 2.340000 0.785000 ;
      RECT 1.875000  0.085000 2.205000 0.445000 ;
      RECT 1.955000  1.835000 2.270000 2.635000 ;
      RECT 1.970000  0.785000 2.340000 1.095000 ;
      RECT 1.970000  1.095000 2.140000 1.495000 ;
      RECT 2.470000  1.355000 2.755000 1.685000 ;
      RECT 2.715000  0.705000 3.095000 1.035000 ;
      RECT 2.745000  2.255000 3.585000 2.425000 ;
      RECT 2.770000  0.365000 3.500000 0.535000 ;
      RECT 2.925000  1.035000 3.095000 1.575000 ;
      RECT 2.925000  1.575000 3.265000 1.905000 ;
      RECT 2.925000  1.905000 3.125000 1.995000 ;
      RECT 3.270000  2.125000 3.585000 2.255000 ;
      RECT 3.305000  2.075000 3.585000 2.125000 ;
      RECT 3.330000  0.535000 3.500000 0.995000 ;
      RECT 3.330000  0.995000 4.200000 1.165000 ;
      RECT 3.395000  2.015000 3.605000 2.045000 ;
      RECT 3.395000  2.045000 3.585000 2.075000 ;
      RECT 3.415000  1.990000 3.605000 2.015000 ;
      RECT 3.420000  1.975000 3.605000 1.990000 ;
      RECT 3.430000  1.960000 3.605000 1.975000 ;
      RECT 3.435000  1.165000 4.200000 1.325000 ;
      RECT 3.435000  1.325000 3.605000 1.960000 ;
      RECT 3.740000  0.085000 4.070000 0.530000 ;
      RECT 3.755000  2.135000 4.600000 2.635000 ;
      RECT 3.840000  1.535000 5.510000 1.705000 ;
      RECT 3.840000  1.705000 4.940000 1.865000 ;
      RECT 4.270000  0.415000 4.570000 0.655000 ;
      RECT 4.270000  0.655000 5.510000 0.825000 ;
      RECT 4.770000  1.865000 4.940000 2.435000 ;
      RECT 5.110000  0.085000 5.490000 0.485000 ;
      RECT 5.110000  1.875000 5.490000 2.635000 ;
      RECT 5.320000  0.825000 5.510000 0.995000 ;
      RECT 5.320000  0.995000 5.620000 1.325000 ;
      RECT 5.320000  1.325000 5.510000 1.535000 ;
      RECT 6.020000  0.085000 6.360000 0.465000 ;
      RECT 6.100000  1.830000 6.360000 2.635000 ;
      RECT 6.535000  0.255000 6.865000 0.995000 ;
      RECT 6.535000  0.995000 7.425000 1.325000 ;
      RECT 6.535000  1.325000 6.870000 2.465000 ;
      RECT 7.035000  0.085000 7.340000 0.545000 ;
      RECT 7.045000  1.835000 7.340000 2.635000 ;
      RECT 7.935000  0.085000 8.195000 0.885000 ;
      RECT 7.935000  1.495000 8.195000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.610000  1.445000 0.780000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.070000  1.785000 1.240000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.470000  1.445000 2.640000 1.615000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 2.930000  1.785000 3.100000 1.955000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
    LAYER met1 ;
      RECT 0.550000 1.415000 0.840000 1.460000 ;
      RECT 0.550000 1.460000 2.700000 1.600000 ;
      RECT 0.550000 1.600000 0.840000 1.645000 ;
      RECT 1.010000 1.755000 1.300000 1.800000 ;
      RECT 1.010000 1.800000 3.160000 1.940000 ;
      RECT 1.010000 1.940000 1.300000 1.985000 ;
      RECT 2.410000 1.415000 2.700000 1.460000 ;
      RECT 2.410000 1.600000 2.700000 1.645000 ;
      RECT 2.870000 1.755000 3.160000 1.800000 ;
      RECT 2.870000 1.940000 3.160000 1.985000 ;
  END
END sky130_fd_sc_hd__dlrbp_2
MACRO sky130_fd_sc_hd__a2bb2oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 0.995000 0.520000 1.615000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.725000 1.010000 1.240000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.780000 0.995000 3.070000 1.615000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.245000 0.995000 2.610000 1.615000 ;
        RECT 2.440000 0.425000 2.610000 0.995000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.515500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 1.785000 1.945000 1.955000 ;
        RECT 1.420000 1.955000 1.785000 2.465000 ;
        RECT 1.775000 0.255000 2.205000 0.825000 ;
        RECT 1.775000 0.825000 1.945000 1.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.220000 0.085000 ;
      RECT 0.000000  2.635000 3.220000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.825000 ;
      RECT 0.095000  1.805000 0.425000 2.635000 ;
      RECT 0.595000  0.255000 0.765000 0.660000 ;
      RECT 0.595000  0.660000 1.580000 0.830000 ;
      RECT 0.875000  1.445000 1.580000 1.615000 ;
      RECT 0.875000  1.615000 1.205000 2.465000 ;
      RECT 0.935000  0.085000 1.605000 0.490000 ;
      RECT 1.410000  0.830000 1.580000 1.445000 ;
      RECT 1.955000  2.235000 2.285000 2.465000 ;
      RECT 2.115000  1.785000 3.130000 1.955000 ;
      RECT 2.115000  1.955000 2.285000 2.235000 ;
      RECT 2.455000  2.135000 2.705000 2.635000 ;
      RECT 2.795000  0.085000 3.125000 0.825000 ;
      RECT 2.875000  1.955000 3.130000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
  END
END sky130_fd_sc_hd__a2bb2oi_1
MACRO sky130_fd_sc_hd__a2bb2oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.945000 1.075000 7.320000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.595000 1.075000 9.045000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 1.555000 1.285000 ;
        RECT 1.385000 1.285000 1.555000 1.445000 ;
        RECT 1.385000 1.445000 3.575000 1.615000 ;
        RECT 3.245000 1.075000 3.575000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.725000 1.075000 3.075000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775000 0.645000 2.995000 0.725000 ;
        RECT 1.775000 0.725000 5.045000 0.905000 ;
        RECT 3.745000 0.905000 3.915000 1.415000 ;
        RECT 3.745000 1.415000 4.965000 1.615000 ;
        RECT 3.875000 0.275000 4.205000 0.725000 ;
        RECT 3.915000 1.615000 4.165000 2.125000 ;
        RECT 4.715000 0.275000 5.045000 0.725000 ;
        RECT 4.745000 1.615000 4.965000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.850000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.085000  1.455000 1.215000 1.625000 ;
      RECT 0.085000  1.625000 0.425000 2.465000 ;
      RECT 0.175000  0.085000 0.345000 0.895000 ;
      RECT 0.515000  0.255000 0.845000 0.725000 ;
      RECT 0.515000  0.725000 1.605000 0.905000 ;
      RECT 0.595000  1.795000 0.805000 2.635000 ;
      RECT 0.975000  1.625000 1.215000 1.795000 ;
      RECT 0.975000  1.795000 3.745000 1.965000 ;
      RECT 0.975000  1.965000 1.215000 2.465000 ;
      RECT 1.015000  0.085000 1.185000 0.555000 ;
      RECT 1.355000  0.255000 3.365000 0.475000 ;
      RECT 1.355000  0.475000 1.605000 0.725000 ;
      RECT 1.395000  2.135000 1.645000 2.635000 ;
      RECT 1.815000  1.965000 2.065000 2.465000 ;
      RECT 2.235000  2.135000 2.485000 2.635000 ;
      RECT 2.655000  1.965000 2.905000 2.465000 ;
      RECT 3.075000  2.135000 3.325000 2.635000 ;
      RECT 3.495000  1.965000 3.745000 2.295000 ;
      RECT 3.495000  2.295000 5.465000 2.465000 ;
      RECT 3.535000  0.085000 3.705000 0.555000 ;
      RECT 4.085000  1.075000 5.725000 1.245000 ;
      RECT 4.335000  1.795000 4.575000 2.295000 ;
      RECT 4.375000  0.085000 4.545000 0.555000 ;
      RECT 5.135000  1.455000 5.465000 2.295000 ;
      RECT 5.215000  0.085000 5.905000 0.555000 ;
      RECT 5.555000  0.735000 9.575000 0.905000 ;
      RECT 5.555000  0.905000 5.725000 1.075000 ;
      RECT 5.655000  1.455000 7.625000 1.625000 ;
      RECT 5.655000  1.625000 5.985000 2.465000 ;
      RECT 6.075000  0.255000 6.405000 0.725000 ;
      RECT 6.075000  0.725000 8.925000 0.735000 ;
      RECT 6.155000  1.795000 6.365000 2.635000 ;
      RECT 6.540000  1.625000 6.780000 2.465000 ;
      RECT 6.575000  0.085000 6.745000 0.555000 ;
      RECT 6.915000  0.255000 7.245000 0.725000 ;
      RECT 6.955000  1.795000 7.205000 2.635000 ;
      RECT 7.375000  1.625000 7.625000 2.295000 ;
      RECT 7.375000  2.295000 9.310000 2.465000 ;
      RECT 7.415000  0.085000 7.585000 0.555000 ;
      RECT 7.755000  0.255000 8.085000 0.725000 ;
      RECT 7.795000  1.455000 9.575000 1.625000 ;
      RECT 7.795000  1.625000 8.045000 2.125000 ;
      RECT 8.215000  1.795000 8.465000 2.295000 ;
      RECT 8.255000  0.085000 8.425000 0.555000 ;
      RECT 8.595000  0.255000 8.925000 0.725000 ;
      RECT 8.635000  1.625000 8.885000 2.125000 ;
      RECT 9.060000  1.795000 9.310000 2.295000 ;
      RECT 9.095000  0.085000 9.265000 0.555000 ;
      RECT 9.215000  0.905000 9.575000 1.455000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
END sky130_fd_sc_hd__a2bb2oi_4
MACRO sky130_fd_sc_hd__a2bb2oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.310000 1.075000 4.205000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.455000 1.075000 5.435000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.710000 1.445000 ;
        RECT 0.085000 1.445000 2.030000 1.615000 ;
        RECT 1.700000 1.075000 2.030000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.940000 1.075000 1.480000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.070000 0.645000 1.400000 0.725000 ;
        RECT 1.070000 0.725000 2.660000 0.905000 ;
        RECT 2.330000 0.255000 2.660000 0.725000 ;
        RECT 2.370000 0.905000 2.660000 1.660000 ;
        RECT 2.370000 1.660000 2.620000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.710000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.520000 0.085000 ;
      RECT 0.000000  2.635000 5.520000 2.805000 ;
      RECT 0.270000  1.785000 2.200000 1.955000 ;
      RECT 0.270000  1.955000 0.520000 2.465000 ;
      RECT 0.310000  0.085000 0.480000 0.895000 ;
      RECT 0.650000  0.255000 1.820000 0.475000 ;
      RECT 0.650000  0.475000 0.900000 0.895000 ;
      RECT 0.690000  2.135000 0.940000 2.635000 ;
      RECT 1.110000  1.955000 1.360000 2.465000 ;
      RECT 1.530000  2.135000 1.780000 2.635000 ;
      RECT 1.950000  1.955000 2.200000 2.295000 ;
      RECT 1.950000  2.295000 3.040000 2.465000 ;
      RECT 1.990000  0.085000 2.160000 0.555000 ;
      RECT 2.790000  1.795000 3.040000 2.295000 ;
      RECT 2.830000  0.085000 3.520000 0.555000 ;
      RECT 2.830000  0.995000 3.120000 1.325000 ;
      RECT 2.950000  0.725000 4.860000 0.905000 ;
      RECT 2.950000  0.905000 3.120000 0.995000 ;
      RECT 2.950000  1.325000 3.120000 1.445000 ;
      RECT 2.950000  1.445000 4.820000 1.615000 ;
      RECT 3.310000  1.785000 4.400000 1.965000 ;
      RECT 3.310000  1.965000 3.560000 2.465000 ;
      RECT 3.690000  0.255000 4.020000 0.725000 ;
      RECT 3.730000  2.135000 3.980000 2.635000 ;
      RECT 4.150000  1.965000 4.400000 2.295000 ;
      RECT 4.150000  2.295000 5.240000 2.465000 ;
      RECT 4.190000  0.085000 4.360000 0.555000 ;
      RECT 4.530000  0.255000 4.860000 0.725000 ;
      RECT 4.570000  1.615000 4.820000 2.125000 ;
      RECT 4.990000  1.455000 5.240000 2.295000 ;
      RECT 5.030000  0.085000 5.200000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
  END
END sky130_fd_sc_hd__a2bb2oi_2
MACRO sky130_fd_sc_hd__clkdlybuf4s18_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s18_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.560000 1.290000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.397600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705000 0.270000 3.150000 0.640000 ;
        RECT 2.715000 1.420000 3.180000 1.525000 ;
        RECT 2.715000 1.525000 3.150000 2.465000 ;
        RECT 2.965000 0.640000 3.150000 0.780000 ;
        RECT 2.965000 0.780000 3.180000 0.945000 ;
        RECT 3.010000 0.945000 3.180000 1.420000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.270000 0.415000 0.735000 ;
      RECT 0.085000  0.735000 1.055000 0.905000 ;
      RECT 0.085000  1.460000 1.055000 1.630000 ;
      RECT 0.085000  1.630000 0.430000 2.465000 ;
      RECT 0.585000  0.085000 0.915000 0.565000 ;
      RECT 0.600000  1.800000 0.930000 2.635000 ;
      RECT 0.730000  0.905000 1.055000 1.460000 ;
      RECT 1.110000  1.800000 1.440000 2.465000 ;
      RECT 1.160000  0.270000 1.440000 0.600000 ;
      RECT 1.270000  0.600000 1.440000 1.075000 ;
      RECT 1.270000  1.075000 2.205000 1.255000 ;
      RECT 1.270000  1.255000 1.440000 1.800000 ;
      RECT 1.630000  0.270000 1.960000 0.735000 ;
      RECT 1.630000  0.735000 2.545000 0.905000 ;
      RECT 1.630000  1.460000 2.545000 1.630000 ;
      RECT 1.630000  1.630000 1.960000 2.465000 ;
      RECT 2.130000  1.800000 2.545000 2.635000 ;
      RECT 2.165000  0.085000 2.535000 0.565000 ;
      RECT 2.375000  0.905000 2.545000 1.075000 ;
      RECT 2.375000  1.075000 2.840000 1.245000 ;
      RECT 2.375000  1.245000 2.545000 1.460000 ;
      RECT 3.320000  0.085000 3.595000 0.645000 ;
      RECT 3.320000  1.625000 3.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s18_2
MACRO sky130_fd_sc_hd__clkdlybuf4s18_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s18_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.055000 0.550000 1.325000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.376300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.210000 0.255000 3.590000 0.545000 ;
        RECT 3.220000 1.760000 3.590000 2.465000 ;
        RECT 3.365000 0.545000 3.590000 1.760000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  0.255000 0.425000 0.715000 ;
      RECT 0.095000  0.715000 1.215000 0.885000 ;
      RECT 0.095000  1.495000 1.215000 1.665000 ;
      RECT 0.095000  1.665000 0.425000 2.465000 ;
      RECT 0.595000  0.085000 0.910000 0.545000 ;
      RECT 0.595000  1.835000 0.925000 2.635000 ;
      RECT 0.720000  0.885000 1.215000 1.495000 ;
      RECT 1.385000  0.255000 1.760000 0.825000 ;
      RECT 1.385000  1.835000 1.760000 2.465000 ;
      RECT 1.590000  0.825000 1.760000 1.055000 ;
      RECT 1.590000  1.055000 2.685000 1.250000 ;
      RECT 1.590000  1.250000 1.760000 1.835000 ;
      RECT 1.930000  0.255000 2.260000 0.715000 ;
      RECT 1.930000  0.715000 3.195000 0.885000 ;
      RECT 1.930000  1.420000 3.195000 1.590000 ;
      RECT 1.930000  1.590000 2.260000 2.465000 ;
      RECT 2.710000  0.085000 3.040000 0.545000 ;
      RECT 2.710000  1.760000 3.040000 2.635000 ;
      RECT 2.855000  0.885000 3.195000 1.420000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s18_1
END LIBRARY