magic
tech sky130A
magscale 1 2
timestamp 1614532237
<< checkpaint >>
rect -3932 -3932 26790 28934
<< viali >>
rect 2053 22049 2087 22083
rect 12817 22049 12851 22083
rect 13921 22049 13955 22083
rect 2237 21845 2271 21879
rect 13001 21845 13035 21879
rect 14105 21845 14139 21879
rect 3617 21641 3651 21675
rect 13645 21641 13679 21675
rect 2605 21437 2639 21471
rect 2697 21437 2731 21471
rect 3157 21437 3191 21471
rect 3341 21437 3375 21471
rect 4629 21437 4663 21471
rect 12633 21437 12667 21471
rect 12725 21437 12759 21471
rect 13093 21437 13127 21471
rect 13185 21437 13219 21471
rect 4813 21301 4847 21335
rect 5273 21097 5307 21131
rect 13185 21097 13219 21131
rect 2053 20961 2087 20995
rect 2421 20961 2455 20995
rect 4077 20961 4111 20995
rect 5181 20961 5215 20995
rect 10885 20961 10919 20995
rect 12173 20961 12207 20995
rect 12725 20961 12759 20995
rect 12909 20961 12943 20995
rect 15301 20961 15335 20995
rect 2145 20893 2179 20927
rect 2329 20893 2363 20927
rect 11989 20893 12023 20927
rect 1685 20825 1719 20859
rect 4261 20757 4295 20791
rect 11069 20757 11103 20791
rect 15485 20757 15519 20791
rect 14657 20553 14691 20587
rect 3801 20485 3835 20519
rect 1501 20417 1535 20451
rect 13001 20417 13035 20451
rect 13369 20417 13403 20451
rect 1593 20349 1627 20383
rect 2053 20349 2087 20383
rect 2145 20349 2179 20383
rect 3617 20349 3651 20383
rect 4721 20349 4755 20383
rect 13093 20349 13127 20383
rect 13461 20349 13495 20383
rect 14473 20349 14507 20383
rect 2605 20213 2639 20247
rect 4905 20213 4939 20247
rect 12725 20213 12759 20247
rect 4261 20009 4295 20043
rect 14013 20009 14047 20043
rect 2237 19941 2271 19975
rect 13001 19941 13035 19975
rect 1777 19873 1811 19907
rect 4077 19873 4111 19907
rect 12449 19873 12483 19907
rect 12541 19873 12575 19907
rect 13829 19873 13863 19907
rect 1685 19805 1719 19839
rect 2053 19261 2087 19295
rect 3157 19261 3191 19295
rect 4261 19261 4295 19295
rect 5365 19261 5399 19295
rect 12817 19261 12851 19295
rect 2237 19125 2271 19159
rect 3341 19125 3375 19159
rect 4445 19125 4479 19159
rect 5549 19125 5583 19159
rect 13001 19125 13035 19159
rect 6469 18921 6503 18955
rect 1685 18785 1719 18819
rect 1777 18785 1811 18819
rect 2237 18785 2271 18819
rect 2421 18785 2455 18819
rect 4077 18785 4111 18819
rect 5181 18785 5215 18819
rect 6285 18785 6319 18819
rect 5365 18649 5399 18683
rect 2697 18581 2731 18615
rect 4261 18581 4295 18615
rect 2145 18377 2179 18411
rect 2329 18241 2363 18275
rect 2513 18173 2547 18207
rect 2881 18173 2915 18207
rect 3065 18173 3099 18207
rect 3893 18173 3927 18207
rect 4445 18173 4479 18207
rect 4721 18173 4755 18207
rect 4905 18173 4939 18207
rect 1409 17697 1443 17731
rect 2605 17697 2639 17731
rect 4077 17697 4111 17731
rect 2513 17629 2547 17663
rect 1593 17493 1627 17527
rect 2789 17493 2823 17527
rect 4261 17493 4295 17527
rect 2881 17289 2915 17323
rect 1777 17221 1811 17255
rect 1685 17085 1719 17119
rect 2697 17085 2731 17119
rect 3801 17085 3835 17119
rect 3985 16949 4019 16983
rect 3065 16745 3099 16779
rect 2881 16609 2915 16643
rect 19717 12733 19751 12767
rect 19901 12597 19935 12631
rect 18337 12257 18371 12291
rect 19533 12257 19567 12291
rect 19441 12189 19475 12223
rect 18521 12053 18555 12087
rect 19717 12053 19751 12087
rect 18153 11645 18187 11679
rect 19441 11645 19475 11679
rect 19533 11645 19567 11679
rect 19993 11645 20027 11679
rect 20177 11645 20211 11679
rect 18337 11509 18371 11543
rect 20453 11509 20487 11543
rect 16773 11305 16807 11339
rect 17877 11305 17911 11339
rect 18797 11237 18831 11271
rect 10793 11169 10827 11203
rect 12357 11169 12391 11203
rect 13461 11169 13495 11203
rect 16589 11169 16623 11203
rect 17693 11169 17727 11203
rect 19441 11169 19475 11203
rect 19809 11169 19843 11203
rect 19993 11169 20027 11203
rect 19533 11101 19567 11135
rect 10977 11033 11011 11067
rect 12541 10965 12575 10999
rect 13645 10965 13679 10999
rect 13829 10761 13863 10795
rect 10517 10625 10551 10659
rect 15761 10625 15795 10659
rect 19349 10625 19383 10659
rect 10425 10557 10459 10591
rect 10793 10557 10827 10591
rect 10885 10557 10919 10591
rect 12817 10557 12851 10591
rect 12909 10557 12943 10591
rect 13277 10557 13311 10591
rect 13369 10557 13403 10591
rect 15301 10557 15335 10591
rect 15485 10557 15519 10591
rect 15853 10557 15887 10591
rect 18153 10557 18187 10591
rect 19441 10557 19475 10591
rect 19993 10557 20027 10591
rect 20177 10557 20211 10591
rect 10057 10421 10091 10455
rect 15117 10421 15151 10455
rect 18337 10421 18371 10455
rect 20453 10421 20487 10455
rect 19073 10217 19107 10251
rect 10609 10149 10643 10183
rect 12817 10149 12851 10183
rect 14381 10149 14415 10183
rect 10149 10081 10183 10115
rect 11529 10081 11563 10115
rect 11713 10081 11747 10115
rect 12265 10081 12299 10115
rect 12449 10081 12483 10115
rect 13921 10081 13955 10115
rect 15301 10081 15335 10115
rect 15485 10081 15519 10115
rect 15945 10081 15979 10115
rect 16037 10081 16071 10115
rect 17693 10081 17727 10115
rect 19441 10081 19475 10115
rect 19809 10081 19843 10115
rect 10057 10013 10091 10047
rect 13829 10013 13863 10047
rect 19533 10013 19567 10047
rect 19717 10013 19751 10047
rect 16405 9945 16439 9979
rect 17877 9877 17911 9911
rect 15117 9537 15151 9571
rect 9873 9469 9907 9503
rect 9965 9469 9999 9503
rect 10425 9469 10459 9503
rect 10609 9469 10643 9503
rect 12449 9469 12483 9503
rect 12541 9469 12575 9503
rect 14013 9469 14047 9503
rect 14105 9469 14139 9503
rect 14473 9469 14507 9503
rect 14565 9469 14599 9503
rect 19441 9469 19475 9503
rect 19533 9469 19567 9503
rect 19991 9469 20025 9503
rect 20177 9469 20211 9503
rect 13001 9401 13035 9435
rect 10885 9333 10919 9367
rect 20453 9333 20487 9367
rect 10793 8993 10827 9027
rect 10885 8993 10919 9027
rect 11345 8993 11379 9027
rect 11529 8993 11563 9027
rect 13277 8993 13311 9027
rect 13461 8993 13495 9027
rect 13829 8993 13863 9027
rect 19533 8993 19567 9027
rect 12817 8925 12851 8959
rect 13737 8925 13771 8959
rect 19441 8925 19475 8959
rect 11805 8789 11839 8823
rect 19717 8789 19751 8823
rect 11437 8585 11471 8619
rect 20361 8517 20395 8551
rect 11253 8381 11287 8415
rect 19441 8381 19475 8415
rect 19533 8381 19567 8415
rect 19901 8381 19935 8415
rect 19993 8381 20027 8415
<< metal1 >>
rect 1104 22330 21712 22352
rect 1104 22278 7851 22330
rect 7903 22278 7915 22330
rect 7967 22278 7979 22330
rect 8031 22278 8043 22330
rect 8095 22278 14720 22330
rect 14772 22278 14784 22330
rect 14836 22278 14848 22330
rect 14900 22278 14912 22330
rect 14964 22278 21712 22330
rect 1104 22256 21712 22278
rect 2041 22083 2099 22089
rect 2041 22049 2053 22083
rect 2087 22080 2099 22083
rect 4246 22080 4252 22092
rect 2087 22052 4252 22080
rect 2087 22049 2099 22052
rect 2041 22043 2099 22049
rect 4246 22040 4252 22052
rect 4304 22040 4310 22092
rect 12805 22083 12863 22089
rect 12805 22049 12817 22083
rect 12851 22049 12863 22083
rect 12805 22043 12863 22049
rect 12820 22012 12848 22043
rect 13170 22040 13176 22092
rect 13228 22080 13234 22092
rect 13909 22083 13967 22089
rect 13909 22080 13921 22083
rect 13228 22052 13921 22080
rect 13228 22040 13234 22052
rect 13909 22049 13921 22052
rect 13955 22049 13967 22083
rect 13909 22043 13967 22049
rect 14550 22012 14556 22024
rect 12820 21984 14556 22012
rect 14550 21972 14556 21984
rect 14608 21972 14614 22024
rect 2225 21879 2283 21885
rect 2225 21845 2237 21879
rect 2271 21876 2283 21879
rect 4706 21876 4712 21888
rect 2271 21848 4712 21876
rect 2271 21845 2283 21848
rect 2225 21839 2283 21845
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 12986 21876 12992 21888
rect 12947 21848 12992 21876
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 13814 21836 13820 21888
rect 13872 21876 13878 21888
rect 14093 21879 14151 21885
rect 14093 21876 14105 21879
rect 13872 21848 14105 21876
rect 13872 21836 13878 21848
rect 14093 21845 14105 21848
rect 14139 21845 14151 21879
rect 14093 21839 14151 21845
rect 1104 21786 21712 21808
rect 1104 21734 4416 21786
rect 4468 21734 4480 21786
rect 4532 21734 4544 21786
rect 4596 21734 4608 21786
rect 4660 21734 11286 21786
rect 11338 21734 11350 21786
rect 11402 21734 11414 21786
rect 11466 21734 11478 21786
rect 11530 21734 18155 21786
rect 18207 21734 18219 21786
rect 18271 21734 18283 21786
rect 18335 21734 18347 21786
rect 18399 21734 21712 21786
rect 1104 21712 21712 21734
rect 3605 21675 3663 21681
rect 3605 21641 3617 21675
rect 3651 21672 3663 21675
rect 4798 21672 4804 21684
rect 3651 21644 4804 21672
rect 3651 21641 3663 21644
rect 3605 21635 3663 21641
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 13446 21632 13452 21684
rect 13504 21672 13510 21684
rect 13633 21675 13691 21681
rect 13633 21672 13645 21675
rect 13504 21644 13645 21672
rect 13504 21632 13510 21644
rect 13633 21641 13645 21644
rect 13679 21641 13691 21675
rect 13633 21635 13691 21641
rect 2608 21508 2820 21536
rect 2608 21477 2636 21508
rect 2593 21471 2651 21477
rect 2593 21437 2605 21471
rect 2639 21437 2651 21471
rect 2593 21431 2651 21437
rect 2685 21471 2743 21477
rect 2685 21437 2697 21471
rect 2731 21437 2743 21471
rect 2792 21468 2820 21508
rect 12636 21508 12848 21536
rect 3142 21468 3148 21480
rect 2792 21440 3148 21468
rect 2685 21431 2743 21437
rect 2700 21400 2728 21431
rect 3142 21428 3148 21440
rect 3200 21428 3206 21480
rect 3326 21468 3332 21480
rect 3287 21440 3332 21468
rect 3326 21428 3332 21440
rect 3384 21428 3390 21480
rect 12636 21477 12664 21508
rect 4617 21471 4675 21477
rect 4617 21468 4629 21471
rect 3436 21440 4629 21468
rect 3344 21400 3372 21428
rect 2700 21372 3372 21400
rect 2038 21292 2044 21344
rect 2096 21332 2102 21344
rect 3436 21332 3464 21440
rect 4617 21437 4629 21440
rect 4663 21437 4675 21471
rect 4617 21431 4675 21437
rect 12621 21471 12679 21477
rect 12621 21437 12633 21471
rect 12667 21437 12679 21471
rect 12621 21431 12679 21437
rect 12713 21471 12771 21477
rect 12713 21437 12725 21471
rect 12759 21437 12771 21471
rect 12820 21468 12848 21508
rect 13078 21468 13084 21480
rect 12820 21440 13084 21468
rect 12713 21431 12771 21437
rect 12728 21400 12756 21431
rect 13078 21428 13084 21440
rect 13136 21428 13142 21480
rect 13173 21471 13231 21477
rect 13173 21437 13185 21471
rect 13219 21437 13231 21471
rect 13173 21431 13231 21437
rect 12986 21400 12992 21412
rect 12728 21372 12992 21400
rect 12986 21360 12992 21372
rect 13044 21400 13050 21412
rect 13188 21400 13216 21431
rect 13044 21372 13216 21400
rect 13044 21360 13050 21372
rect 14090 21360 14096 21412
rect 14148 21400 14154 21412
rect 19334 21400 19340 21412
rect 14148 21372 19340 21400
rect 14148 21360 14154 21372
rect 19334 21360 19340 21372
rect 19392 21360 19398 21412
rect 2096 21304 3464 21332
rect 2096 21292 2102 21304
rect 4062 21292 4068 21344
rect 4120 21332 4126 21344
rect 4801 21335 4859 21341
rect 4801 21332 4813 21335
rect 4120 21304 4813 21332
rect 4120 21292 4126 21304
rect 4801 21301 4813 21304
rect 4847 21301 4859 21335
rect 4801 21295 4859 21301
rect 1104 21242 21712 21264
rect 1104 21190 7851 21242
rect 7903 21190 7915 21242
rect 7967 21190 7979 21242
rect 8031 21190 8043 21242
rect 8095 21190 14720 21242
rect 14772 21190 14784 21242
rect 14836 21190 14848 21242
rect 14900 21190 14912 21242
rect 14964 21190 21712 21242
rect 1104 21168 21712 21190
rect 2222 21088 2228 21140
rect 2280 21128 2286 21140
rect 2280 21100 3280 21128
rect 2280 21088 2286 21100
rect 1578 21020 1584 21072
rect 1636 21060 1642 21072
rect 3252 21060 3280 21100
rect 3326 21088 3332 21140
rect 3384 21128 3390 21140
rect 5261 21131 5319 21137
rect 5261 21128 5273 21131
rect 3384 21100 5273 21128
rect 3384 21088 3390 21100
rect 5261 21097 5273 21100
rect 5307 21097 5319 21131
rect 5261 21091 5319 21097
rect 13078 21088 13084 21140
rect 13136 21128 13142 21140
rect 13173 21131 13231 21137
rect 13173 21128 13185 21131
rect 13136 21100 13185 21128
rect 13136 21088 13142 21100
rect 13173 21097 13185 21100
rect 13219 21097 13231 21131
rect 13173 21091 13231 21097
rect 12434 21060 12440 21072
rect 1636 21032 2452 21060
rect 3252 21032 5212 21060
rect 1636 21020 1642 21032
rect 2038 20992 2044 21004
rect 1999 20964 2044 20992
rect 2038 20952 2044 20964
rect 2096 20952 2102 21004
rect 2424 21001 2452 21032
rect 2409 20995 2467 21001
rect 2409 20961 2421 20995
rect 2455 20961 2467 20995
rect 4062 20992 4068 21004
rect 4023 20964 4068 20992
rect 2409 20955 2467 20961
rect 4062 20952 4068 20964
rect 4120 20952 4126 21004
rect 5184 21001 5212 21032
rect 11992 21032 12440 21060
rect 5169 20995 5227 21001
rect 5169 20961 5181 20995
rect 5215 20961 5227 20995
rect 5169 20955 5227 20961
rect 10873 20995 10931 21001
rect 10873 20961 10885 20995
rect 10919 20992 10931 20995
rect 11882 20992 11888 21004
rect 10919 20964 11888 20992
rect 10919 20961 10931 20964
rect 10873 20955 10931 20961
rect 11882 20952 11888 20964
rect 11940 20952 11946 21004
rect 2130 20924 2136 20936
rect 2091 20896 2136 20924
rect 2130 20884 2136 20896
rect 2188 20884 2194 20936
rect 2314 20924 2320 20936
rect 2275 20896 2320 20924
rect 2314 20884 2320 20896
rect 2372 20884 2378 20936
rect 7742 20884 7748 20936
rect 7800 20924 7806 20936
rect 11992 20933 12020 21032
rect 12434 21020 12440 21032
rect 12492 21060 12498 21072
rect 12492 21032 12940 21060
rect 12492 21020 12498 21032
rect 12161 20995 12219 21001
rect 12161 20961 12173 20995
rect 12207 20992 12219 20995
rect 12710 20992 12716 21004
rect 12207 20964 12716 20992
rect 12207 20961 12219 20964
rect 12161 20955 12219 20961
rect 12710 20952 12716 20964
rect 12768 20952 12774 21004
rect 12912 21001 12940 21032
rect 12897 20995 12955 21001
rect 12897 20961 12909 20995
rect 12943 20992 12955 20995
rect 13354 20992 13360 21004
rect 12943 20964 13360 20992
rect 12943 20961 12955 20964
rect 12897 20955 12955 20961
rect 13354 20952 13360 20964
rect 13412 20952 13418 21004
rect 15286 20992 15292 21004
rect 15247 20964 15292 20992
rect 15286 20952 15292 20964
rect 15344 20952 15350 21004
rect 11977 20927 12035 20933
rect 11977 20924 11989 20927
rect 7800 20896 11989 20924
rect 7800 20884 7806 20896
rect 11977 20893 11989 20896
rect 12023 20893 12035 20927
rect 11977 20887 12035 20893
rect 1673 20859 1731 20865
rect 1673 20825 1685 20859
rect 1719 20856 1731 20859
rect 13078 20856 13084 20868
rect 1719 20828 13084 20856
rect 1719 20825 1731 20828
rect 1673 20819 1731 20825
rect 13078 20816 13084 20828
rect 13136 20816 13142 20868
rect 4246 20788 4252 20800
rect 4207 20760 4252 20788
rect 4246 20748 4252 20760
rect 4304 20748 4310 20800
rect 11057 20791 11115 20797
rect 11057 20757 11069 20791
rect 11103 20788 11115 20791
rect 12802 20788 12808 20800
rect 11103 20760 12808 20788
rect 11103 20757 11115 20760
rect 11057 20751 11115 20757
rect 12802 20748 12808 20760
rect 12860 20748 12866 20800
rect 15470 20788 15476 20800
rect 15431 20760 15476 20788
rect 15470 20748 15476 20760
rect 15528 20748 15534 20800
rect 1104 20698 21712 20720
rect 1104 20646 4416 20698
rect 4468 20646 4480 20698
rect 4532 20646 4544 20698
rect 4596 20646 4608 20698
rect 4660 20646 11286 20698
rect 11338 20646 11350 20698
rect 11402 20646 11414 20698
rect 11466 20646 11478 20698
rect 11530 20646 18155 20698
rect 18207 20646 18219 20698
rect 18271 20646 18283 20698
rect 18335 20646 18347 20698
rect 18399 20646 21712 20698
rect 1104 20624 21712 20646
rect 12710 20544 12716 20596
rect 12768 20584 12774 20596
rect 12768 20556 13584 20584
rect 12768 20544 12774 20556
rect 2314 20516 2320 20528
rect 1780 20488 2320 20516
rect 1486 20448 1492 20460
rect 1447 20420 1492 20448
rect 1486 20408 1492 20420
rect 1544 20448 1550 20460
rect 1780 20448 1808 20488
rect 2314 20476 2320 20488
rect 2372 20476 2378 20528
rect 3789 20519 3847 20525
rect 3789 20485 3801 20519
rect 3835 20516 3847 20519
rect 4246 20516 4252 20528
rect 3835 20488 4252 20516
rect 3835 20485 3847 20488
rect 3789 20479 3847 20485
rect 4246 20476 4252 20488
rect 4304 20476 4310 20528
rect 13556 20516 13584 20556
rect 14550 20544 14556 20596
rect 14608 20584 14614 20596
rect 14645 20587 14703 20593
rect 14645 20584 14657 20587
rect 14608 20556 14657 20584
rect 14608 20544 14614 20556
rect 14645 20553 14657 20556
rect 14691 20553 14703 20587
rect 14645 20547 14703 20553
rect 13556 20488 16528 20516
rect 12986 20448 12992 20460
rect 1544 20420 1808 20448
rect 12947 20420 12992 20448
rect 1544 20408 1550 20420
rect 1578 20380 1584 20392
rect 1539 20352 1584 20380
rect 1578 20340 1584 20352
rect 1636 20340 1642 20392
rect 1780 20380 1808 20420
rect 12986 20408 12992 20420
rect 13044 20408 13050 20460
rect 13354 20448 13360 20460
rect 13315 20420 13360 20448
rect 13354 20408 13360 20420
rect 13412 20408 13418 20460
rect 2041 20383 2099 20389
rect 2041 20380 2053 20383
rect 1780 20352 2053 20380
rect 2041 20349 2053 20352
rect 2087 20349 2099 20383
rect 2041 20343 2099 20349
rect 2133 20383 2191 20389
rect 2133 20349 2145 20383
rect 2179 20349 2191 20383
rect 3602 20380 3608 20392
rect 3563 20352 3608 20380
rect 2133 20343 2191 20349
rect 1596 20312 1624 20340
rect 2148 20312 2176 20343
rect 3602 20340 3608 20352
rect 3660 20340 3666 20392
rect 4706 20380 4712 20392
rect 4667 20352 4712 20380
rect 4706 20340 4712 20352
rect 4764 20340 4770 20392
rect 13078 20380 13084 20392
rect 13039 20352 13084 20380
rect 13078 20340 13084 20352
rect 13136 20340 13142 20392
rect 13449 20383 13507 20389
rect 13449 20349 13461 20383
rect 13495 20380 13507 20383
rect 13556 20380 13584 20488
rect 15194 20408 15200 20460
rect 15252 20448 15258 20460
rect 16390 20448 16396 20460
rect 15252 20420 16396 20448
rect 15252 20408 15258 20420
rect 16390 20408 16396 20420
rect 16448 20408 16454 20460
rect 16500 20448 16528 20488
rect 18414 20448 18420 20460
rect 16500 20420 18420 20448
rect 18414 20408 18420 20420
rect 18472 20408 18478 20460
rect 20714 20408 20720 20460
rect 20772 20448 20778 20460
rect 22094 20448 22100 20460
rect 20772 20420 22100 20448
rect 20772 20408 20778 20420
rect 22094 20408 22100 20420
rect 22152 20408 22158 20460
rect 13495 20352 13584 20380
rect 14461 20383 14519 20389
rect 13495 20349 13507 20352
rect 13449 20343 13507 20349
rect 14461 20349 14473 20383
rect 14507 20380 14519 20383
rect 15470 20380 15476 20392
rect 14507 20352 15476 20380
rect 14507 20349 14519 20352
rect 14461 20343 14519 20349
rect 15470 20340 15476 20352
rect 15528 20340 15534 20392
rect 1596 20284 2176 20312
rect 2590 20244 2596 20256
rect 2551 20216 2596 20244
rect 2590 20204 2596 20216
rect 2648 20204 2654 20256
rect 4062 20204 4068 20256
rect 4120 20244 4126 20256
rect 4893 20247 4951 20253
rect 4893 20244 4905 20247
rect 4120 20216 4905 20244
rect 4120 20204 4126 20216
rect 4893 20213 4905 20216
rect 4939 20213 4951 20247
rect 4893 20207 4951 20213
rect 12713 20247 12771 20253
rect 12713 20213 12725 20247
rect 12759 20244 12771 20247
rect 17678 20244 17684 20256
rect 12759 20216 17684 20244
rect 12759 20213 12771 20216
rect 12713 20207 12771 20213
rect 17678 20204 17684 20216
rect 17736 20204 17742 20256
rect 1104 20154 21712 20176
rect 1104 20102 7851 20154
rect 7903 20102 7915 20154
rect 7967 20102 7979 20154
rect 8031 20102 8043 20154
rect 8095 20102 14720 20154
rect 14772 20102 14784 20154
rect 14836 20102 14848 20154
rect 14900 20102 14912 20154
rect 14964 20102 21712 20154
rect 1104 20080 21712 20102
rect 3602 20000 3608 20052
rect 3660 20040 3666 20052
rect 4249 20043 4307 20049
rect 4249 20040 4261 20043
rect 3660 20012 4261 20040
rect 3660 20000 3666 20012
rect 4249 20009 4261 20012
rect 4295 20009 4307 20043
rect 4249 20003 4307 20009
rect 11882 20000 11888 20052
rect 11940 20040 11946 20052
rect 14001 20043 14059 20049
rect 14001 20040 14013 20043
rect 11940 20012 14013 20040
rect 11940 20000 11946 20012
rect 14001 20009 14013 20012
rect 14047 20009 14059 20043
rect 14001 20003 14059 20009
rect 2130 19932 2136 19984
rect 2188 19972 2194 19984
rect 2225 19975 2283 19981
rect 2225 19972 2237 19975
rect 2188 19944 2237 19972
rect 2188 19932 2194 19944
rect 2225 19941 2237 19944
rect 2271 19941 2283 19975
rect 12986 19972 12992 19984
rect 12947 19944 12992 19972
rect 2225 19935 2283 19941
rect 12986 19932 12992 19944
rect 13044 19932 13050 19984
rect 1578 19864 1584 19916
rect 1636 19904 1642 19916
rect 1765 19907 1823 19913
rect 1765 19904 1777 19907
rect 1636 19876 1777 19904
rect 1636 19864 1642 19876
rect 1765 19873 1777 19876
rect 1811 19873 1823 19907
rect 4062 19904 4068 19916
rect 4023 19876 4068 19904
rect 1765 19867 1823 19873
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 12434 19904 12440 19916
rect 12395 19876 12440 19904
rect 12434 19864 12440 19876
rect 12492 19864 12498 19916
rect 12529 19907 12587 19913
rect 12529 19873 12541 19907
rect 12575 19904 12587 19907
rect 12710 19904 12716 19916
rect 12575 19876 12716 19904
rect 12575 19873 12587 19876
rect 12529 19867 12587 19873
rect 12710 19864 12716 19876
rect 12768 19864 12774 19916
rect 13814 19904 13820 19916
rect 13775 19876 13820 19904
rect 13814 19864 13820 19876
rect 13872 19864 13878 19916
rect 1486 19796 1492 19848
rect 1544 19836 1550 19848
rect 1673 19839 1731 19845
rect 1673 19836 1685 19839
rect 1544 19808 1685 19836
rect 1544 19796 1550 19808
rect 1673 19805 1685 19808
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 1104 19610 21712 19632
rect 1104 19558 4416 19610
rect 4468 19558 4480 19610
rect 4532 19558 4544 19610
rect 4596 19558 4608 19610
rect 4660 19558 11286 19610
rect 11338 19558 11350 19610
rect 11402 19558 11414 19610
rect 11466 19558 11478 19610
rect 11530 19558 18155 19610
rect 18207 19558 18219 19610
rect 18271 19558 18283 19610
rect 18335 19558 18347 19610
rect 18399 19558 21712 19610
rect 1104 19536 21712 19558
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19292 2099 19295
rect 3145 19295 3203 19301
rect 3145 19292 3157 19295
rect 2087 19264 3157 19292
rect 2087 19261 2099 19264
rect 2041 19255 2099 19261
rect 3145 19261 3157 19264
rect 3191 19261 3203 19295
rect 4246 19292 4252 19304
rect 4207 19264 4252 19292
rect 3145 19255 3203 19261
rect 3160 19224 3188 19255
rect 4246 19252 4252 19264
rect 4304 19252 4310 19304
rect 5353 19295 5411 19301
rect 5353 19261 5365 19295
rect 5399 19292 5411 19295
rect 6454 19292 6460 19304
rect 5399 19264 6460 19292
rect 5399 19261 5411 19264
rect 5353 19255 5411 19261
rect 6454 19252 6460 19264
rect 6512 19252 6518 19304
rect 12802 19292 12808 19304
rect 12763 19264 12808 19292
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 3160 19196 4476 19224
rect 1762 19116 1768 19168
rect 1820 19156 1826 19168
rect 2225 19159 2283 19165
rect 2225 19156 2237 19159
rect 1820 19128 2237 19156
rect 1820 19116 1826 19128
rect 2225 19125 2237 19128
rect 2271 19125 2283 19159
rect 2225 19119 2283 19125
rect 2314 19116 2320 19168
rect 2372 19156 2378 19168
rect 4448 19165 4476 19196
rect 3329 19159 3387 19165
rect 3329 19156 3341 19159
rect 2372 19128 3341 19156
rect 2372 19116 2378 19128
rect 3329 19125 3341 19128
rect 3375 19125 3387 19159
rect 3329 19119 3387 19125
rect 4433 19159 4491 19165
rect 4433 19125 4445 19159
rect 4479 19125 4491 19159
rect 4433 19119 4491 19125
rect 4706 19116 4712 19168
rect 4764 19156 4770 19168
rect 5537 19159 5595 19165
rect 5537 19156 5549 19159
rect 4764 19128 5549 19156
rect 4764 19116 4770 19128
rect 5537 19125 5549 19128
rect 5583 19125 5595 19159
rect 5537 19119 5595 19125
rect 12989 19159 13047 19165
rect 12989 19125 13001 19159
rect 13035 19156 13047 19159
rect 15286 19156 15292 19168
rect 13035 19128 15292 19156
rect 13035 19125 13047 19128
rect 12989 19119 13047 19125
rect 15286 19116 15292 19128
rect 15344 19116 15350 19168
rect 1104 19066 21712 19088
rect 1104 19014 7851 19066
rect 7903 19014 7915 19066
rect 7967 19014 7979 19066
rect 8031 19014 8043 19066
rect 8095 19014 14720 19066
rect 14772 19014 14784 19066
rect 14836 19014 14848 19066
rect 14900 19014 14912 19066
rect 14964 19014 21712 19066
rect 1104 18992 21712 19014
rect 6454 18952 6460 18964
rect 6415 18924 6460 18952
rect 6454 18912 6460 18924
rect 6512 18912 6518 18964
rect 1688 18856 2452 18884
rect 1688 18825 1716 18856
rect 1673 18819 1731 18825
rect 1673 18785 1685 18819
rect 1719 18785 1731 18819
rect 1673 18779 1731 18785
rect 1762 18776 1768 18828
rect 1820 18816 1826 18828
rect 2225 18819 2283 18825
rect 1820 18788 1865 18816
rect 1820 18776 1826 18788
rect 2225 18785 2237 18819
rect 2271 18816 2283 18819
rect 2314 18816 2320 18828
rect 2271 18788 2320 18816
rect 2271 18785 2283 18788
rect 2225 18779 2283 18785
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 2424 18825 2452 18856
rect 2409 18819 2467 18825
rect 2409 18785 2421 18819
rect 2455 18816 2467 18819
rect 2590 18816 2596 18828
rect 2455 18788 2596 18816
rect 2455 18785 2467 18788
rect 2409 18779 2467 18785
rect 2590 18776 2596 18788
rect 2648 18776 2654 18828
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18785 4123 18819
rect 5166 18816 5172 18828
rect 5127 18788 5172 18816
rect 4065 18779 4123 18785
rect 4080 18748 4108 18779
rect 5166 18776 5172 18788
rect 5224 18776 5230 18828
rect 5258 18776 5264 18828
rect 5316 18816 5322 18828
rect 6273 18819 6331 18825
rect 6273 18816 6285 18819
rect 5316 18788 6285 18816
rect 5316 18776 5322 18788
rect 6273 18785 6285 18788
rect 6319 18785 6331 18819
rect 6273 18779 6331 18785
rect 4080 18720 5396 18748
rect 5368 18689 5396 18720
rect 5353 18683 5411 18689
rect 5353 18649 5365 18683
rect 5399 18649 5411 18683
rect 5353 18643 5411 18649
rect 2682 18612 2688 18624
rect 2643 18584 2688 18612
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 4246 18612 4252 18624
rect 4207 18584 4252 18612
rect 4246 18572 4252 18584
rect 4304 18572 4310 18624
rect 1104 18522 21712 18544
rect 1104 18470 4416 18522
rect 4468 18470 4480 18522
rect 4532 18470 4544 18522
rect 4596 18470 4608 18522
rect 4660 18470 11286 18522
rect 11338 18470 11350 18522
rect 11402 18470 11414 18522
rect 11466 18470 11478 18522
rect 11530 18470 18155 18522
rect 18207 18470 18219 18522
rect 18271 18470 18283 18522
rect 18335 18470 18347 18522
rect 18399 18470 21712 18522
rect 1104 18448 21712 18470
rect 2038 18368 2044 18420
rect 2096 18408 2102 18420
rect 2133 18411 2191 18417
rect 2133 18408 2145 18411
rect 2096 18380 2145 18408
rect 2096 18368 2102 18380
rect 2133 18377 2145 18380
rect 2179 18377 2191 18411
rect 2133 18371 2191 18377
rect 2222 18232 2228 18284
rect 2280 18272 2286 18284
rect 2317 18275 2375 18281
rect 2317 18272 2329 18275
rect 2280 18244 2329 18272
rect 2280 18232 2286 18244
rect 2317 18241 2329 18244
rect 2363 18241 2375 18275
rect 2317 18235 2375 18241
rect 2884 18244 4752 18272
rect 2498 18204 2504 18216
rect 2459 18176 2504 18204
rect 2498 18164 2504 18176
rect 2556 18164 2562 18216
rect 2774 18164 2780 18216
rect 2832 18204 2838 18216
rect 2884 18213 2912 18244
rect 2869 18207 2927 18213
rect 2869 18204 2881 18207
rect 2832 18176 2881 18204
rect 2832 18164 2838 18176
rect 2869 18173 2881 18176
rect 2915 18173 2927 18207
rect 3050 18204 3056 18216
rect 2963 18176 3056 18204
rect 2869 18167 2927 18173
rect 3050 18164 3056 18176
rect 3108 18164 3114 18216
rect 3142 18164 3148 18216
rect 3200 18204 3206 18216
rect 3881 18207 3939 18213
rect 3881 18204 3893 18207
rect 3200 18176 3893 18204
rect 3200 18164 3206 18176
rect 3881 18173 3893 18176
rect 3927 18173 3939 18207
rect 3881 18167 3939 18173
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 4724 18213 4752 18244
rect 4433 18207 4491 18213
rect 4433 18204 4445 18207
rect 4212 18176 4445 18204
rect 4212 18164 4218 18176
rect 4433 18173 4445 18176
rect 4479 18173 4491 18207
rect 4433 18167 4491 18173
rect 4709 18207 4767 18213
rect 4709 18173 4721 18207
rect 4755 18173 4767 18207
rect 4709 18167 4767 18173
rect 4893 18207 4951 18213
rect 4893 18173 4905 18207
rect 4939 18173 4951 18207
rect 4893 18167 4951 18173
rect 3068 18136 3096 18164
rect 4908 18136 4936 18167
rect 3068 18108 4936 18136
rect 1104 17978 21712 18000
rect 1104 17926 7851 17978
rect 7903 17926 7915 17978
rect 7967 17926 7979 17978
rect 8031 17926 8043 17978
rect 8095 17926 14720 17978
rect 14772 17926 14784 17978
rect 14836 17926 14848 17978
rect 14900 17926 14912 17978
rect 14964 17926 21712 17978
rect 1104 17904 21712 17926
rect 2498 17796 2504 17808
rect 1412 17768 2504 17796
rect 1412 17737 1440 17768
rect 2498 17756 2504 17768
rect 2556 17756 2562 17808
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17697 1455 17731
rect 1397 17691 1455 17697
rect 2593 17731 2651 17737
rect 2593 17697 2605 17731
rect 2639 17728 2651 17731
rect 2774 17728 2780 17740
rect 2639 17700 2780 17728
rect 2639 17697 2651 17700
rect 2593 17691 2651 17697
rect 2774 17688 2780 17700
rect 2832 17688 2838 17740
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17728 4123 17731
rect 4706 17728 4712 17740
rect 4111 17700 4712 17728
rect 4111 17697 4123 17700
rect 4065 17691 4123 17697
rect 4706 17688 4712 17700
rect 4764 17688 4770 17740
rect 2501 17663 2559 17669
rect 2501 17629 2513 17663
rect 2547 17660 2559 17663
rect 2866 17660 2872 17672
rect 2547 17632 2872 17660
rect 2547 17629 2559 17632
rect 2501 17623 2559 17629
rect 2866 17620 2872 17632
rect 2924 17660 2930 17672
rect 3050 17660 3056 17672
rect 2924 17632 3056 17660
rect 2924 17620 2930 17632
rect 3050 17620 3056 17632
rect 3108 17620 3114 17672
rect 1578 17524 1584 17536
rect 1539 17496 1584 17524
rect 1578 17484 1584 17496
rect 1636 17484 1642 17536
rect 2498 17484 2504 17536
rect 2556 17524 2562 17536
rect 2777 17527 2835 17533
rect 2777 17524 2789 17527
rect 2556 17496 2789 17524
rect 2556 17484 2562 17496
rect 2777 17493 2789 17496
rect 2823 17493 2835 17527
rect 2777 17487 2835 17493
rect 2866 17484 2872 17536
rect 2924 17524 2930 17536
rect 4249 17527 4307 17533
rect 4249 17524 4261 17527
rect 2924 17496 4261 17524
rect 2924 17484 2930 17496
rect 4249 17493 4261 17496
rect 4295 17493 4307 17527
rect 4249 17487 4307 17493
rect 1104 17434 21712 17456
rect 1104 17382 4416 17434
rect 4468 17382 4480 17434
rect 4532 17382 4544 17434
rect 4596 17382 4608 17434
rect 4660 17382 11286 17434
rect 11338 17382 11350 17434
rect 11402 17382 11414 17434
rect 11466 17382 11478 17434
rect 11530 17382 18155 17434
rect 18207 17382 18219 17434
rect 18271 17382 18283 17434
rect 18335 17382 18347 17434
rect 18399 17382 21712 17434
rect 1104 17360 21712 17382
rect 2869 17323 2927 17329
rect 2869 17289 2881 17323
rect 2915 17320 2927 17323
rect 5166 17320 5172 17332
rect 2915 17292 5172 17320
rect 2915 17289 2927 17292
rect 2869 17283 2927 17289
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 1765 17255 1823 17261
rect 1765 17221 1777 17255
rect 1811 17252 1823 17255
rect 4154 17252 4160 17264
rect 1811 17224 4160 17252
rect 1811 17221 1823 17224
rect 1765 17215 1823 17221
rect 4154 17212 4160 17224
rect 4212 17212 4218 17264
rect 1578 17144 1584 17196
rect 1636 17184 1642 17196
rect 1636 17156 3832 17184
rect 1636 17144 1642 17156
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17085 1731 17119
rect 1673 17079 1731 17085
rect 2685 17119 2743 17125
rect 2685 17085 2697 17119
rect 2731 17116 2743 17119
rect 2866 17116 2872 17128
rect 2731 17088 2872 17116
rect 2731 17085 2743 17088
rect 2685 17079 2743 17085
rect 1688 17048 1716 17079
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 3804 17125 3832 17156
rect 3789 17119 3847 17125
rect 3789 17085 3801 17119
rect 3835 17085 3847 17119
rect 3789 17079 3847 17085
rect 4246 17048 4252 17060
rect 1688 17020 4252 17048
rect 4246 17008 4252 17020
rect 4304 17008 4310 17060
rect 3970 16980 3976 16992
rect 3931 16952 3976 16980
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 1104 16890 21712 16912
rect 1104 16838 7851 16890
rect 7903 16838 7915 16890
rect 7967 16838 7979 16890
rect 8031 16838 8043 16890
rect 8095 16838 14720 16890
rect 14772 16838 14784 16890
rect 14836 16838 14848 16890
rect 14900 16838 14912 16890
rect 14964 16838 21712 16890
rect 1104 16816 21712 16838
rect 3053 16779 3111 16785
rect 3053 16745 3065 16779
rect 3099 16776 3111 16779
rect 5258 16776 5264 16788
rect 3099 16748 5264 16776
rect 3099 16745 3111 16748
rect 3053 16739 3111 16745
rect 5258 16736 5264 16748
rect 5316 16736 5322 16788
rect 2869 16643 2927 16649
rect 2869 16609 2881 16643
rect 2915 16640 2927 16643
rect 3970 16640 3976 16652
rect 2915 16612 3976 16640
rect 2915 16609 2927 16612
rect 2869 16603 2927 16609
rect 3970 16600 3976 16612
rect 4028 16600 4034 16652
rect 1104 16346 21712 16368
rect 1104 16294 4416 16346
rect 4468 16294 4480 16346
rect 4532 16294 4544 16346
rect 4596 16294 4608 16346
rect 4660 16294 11286 16346
rect 11338 16294 11350 16346
rect 11402 16294 11414 16346
rect 11466 16294 11478 16346
rect 11530 16294 18155 16346
rect 18207 16294 18219 16346
rect 18271 16294 18283 16346
rect 18335 16294 18347 16346
rect 18399 16294 21712 16346
rect 1104 16272 21712 16294
rect 1104 15802 21712 15824
rect 1104 15750 7851 15802
rect 7903 15750 7915 15802
rect 7967 15750 7979 15802
rect 8031 15750 8043 15802
rect 8095 15750 14720 15802
rect 14772 15750 14784 15802
rect 14836 15750 14848 15802
rect 14900 15750 14912 15802
rect 14964 15750 21712 15802
rect 1104 15728 21712 15750
rect 1104 15258 21712 15280
rect 1104 15206 4416 15258
rect 4468 15206 4480 15258
rect 4532 15206 4544 15258
rect 4596 15206 4608 15258
rect 4660 15206 11286 15258
rect 11338 15206 11350 15258
rect 11402 15206 11414 15258
rect 11466 15206 11478 15258
rect 11530 15206 18155 15258
rect 18207 15206 18219 15258
rect 18271 15206 18283 15258
rect 18335 15206 18347 15258
rect 18399 15206 21712 15258
rect 1104 15184 21712 15206
rect 1104 14714 21712 14736
rect 1104 14662 7851 14714
rect 7903 14662 7915 14714
rect 7967 14662 7979 14714
rect 8031 14662 8043 14714
rect 8095 14662 14720 14714
rect 14772 14662 14784 14714
rect 14836 14662 14848 14714
rect 14900 14662 14912 14714
rect 14964 14662 21712 14714
rect 1104 14640 21712 14662
rect 1104 14170 21712 14192
rect 1104 14118 4416 14170
rect 4468 14118 4480 14170
rect 4532 14118 4544 14170
rect 4596 14118 4608 14170
rect 4660 14118 11286 14170
rect 11338 14118 11350 14170
rect 11402 14118 11414 14170
rect 11466 14118 11478 14170
rect 11530 14118 18155 14170
rect 18207 14118 18219 14170
rect 18271 14118 18283 14170
rect 18335 14118 18347 14170
rect 18399 14118 21712 14170
rect 1104 14096 21712 14118
rect 1104 13626 21712 13648
rect 1104 13574 7851 13626
rect 7903 13574 7915 13626
rect 7967 13574 7979 13626
rect 8031 13574 8043 13626
rect 8095 13574 14720 13626
rect 14772 13574 14784 13626
rect 14836 13574 14848 13626
rect 14900 13574 14912 13626
rect 14964 13574 21712 13626
rect 1104 13552 21712 13574
rect 1104 13082 21712 13104
rect 1104 13030 4416 13082
rect 4468 13030 4480 13082
rect 4532 13030 4544 13082
rect 4596 13030 4608 13082
rect 4660 13030 11286 13082
rect 11338 13030 11350 13082
rect 11402 13030 11414 13082
rect 11466 13030 11478 13082
rect 11530 13030 18155 13082
rect 18207 13030 18219 13082
rect 18271 13030 18283 13082
rect 18335 13030 18347 13082
rect 18399 13030 21712 13082
rect 1104 13008 21712 13030
rect 19334 12724 19340 12776
rect 19392 12764 19398 12776
rect 19705 12767 19763 12773
rect 19705 12764 19717 12767
rect 19392 12736 19717 12764
rect 19392 12724 19398 12736
rect 19705 12733 19717 12736
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 3418 12588 3424 12640
rect 3476 12628 3482 12640
rect 13906 12628 13912 12640
rect 3476 12600 13912 12628
rect 3476 12588 3482 12600
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 19889 12631 19947 12637
rect 19889 12628 19901 12631
rect 19484 12600 19901 12628
rect 19484 12588 19490 12600
rect 19889 12597 19901 12600
rect 19935 12597 19947 12631
rect 19889 12591 19947 12597
rect 1104 12538 21712 12560
rect 1104 12486 7851 12538
rect 7903 12486 7915 12538
rect 7967 12486 7979 12538
rect 8031 12486 8043 12538
rect 8095 12486 14720 12538
rect 14772 12486 14784 12538
rect 14836 12486 14848 12538
rect 14900 12486 14912 12538
rect 14964 12486 21712 12538
rect 1104 12464 21712 12486
rect 16758 12248 16764 12300
rect 16816 12288 16822 12300
rect 18325 12291 18383 12297
rect 18325 12288 18337 12291
rect 16816 12260 18337 12288
rect 16816 12248 16822 12260
rect 18325 12257 18337 12260
rect 18371 12257 18383 12291
rect 19518 12288 19524 12300
rect 19479 12260 19524 12288
rect 18325 12251 18383 12257
rect 19518 12248 19524 12260
rect 19576 12248 19582 12300
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12220 19487 12223
rect 20714 12220 20720 12232
rect 19475 12192 20720 12220
rect 19475 12189 19487 12192
rect 19429 12183 19487 12189
rect 20714 12180 20720 12192
rect 20772 12180 20778 12232
rect 17678 12044 17684 12096
rect 17736 12084 17742 12096
rect 18509 12087 18567 12093
rect 18509 12084 18521 12087
rect 17736 12056 18521 12084
rect 17736 12044 17742 12056
rect 18509 12053 18521 12056
rect 18555 12053 18567 12087
rect 18509 12047 18567 12053
rect 19518 12044 19524 12096
rect 19576 12084 19582 12096
rect 19705 12087 19763 12093
rect 19705 12084 19717 12087
rect 19576 12056 19717 12084
rect 19576 12044 19582 12056
rect 19705 12053 19717 12056
rect 19751 12053 19763 12087
rect 19705 12047 19763 12053
rect 1104 11994 21712 12016
rect 1104 11942 4416 11994
rect 4468 11942 4480 11994
rect 4532 11942 4544 11994
rect 4596 11942 4608 11994
rect 4660 11942 11286 11994
rect 11338 11942 11350 11994
rect 11402 11942 11414 11994
rect 11466 11942 11478 11994
rect 11530 11942 18155 11994
rect 18207 11942 18219 11994
rect 18271 11942 18283 11994
rect 18335 11942 18347 11994
rect 18399 11942 21712 11994
rect 1104 11920 21712 11942
rect 19444 11716 19656 11744
rect 17862 11636 17868 11688
rect 17920 11676 17926 11688
rect 19444 11685 19472 11716
rect 19628 11688 19656 11716
rect 18141 11679 18199 11685
rect 18141 11676 18153 11679
rect 17920 11648 18153 11676
rect 17920 11636 17926 11648
rect 18141 11645 18153 11648
rect 18187 11645 18199 11679
rect 18141 11639 18199 11645
rect 19429 11679 19487 11685
rect 19429 11645 19441 11679
rect 19475 11645 19487 11679
rect 19429 11639 19487 11645
rect 19521 11679 19579 11685
rect 19521 11645 19533 11679
rect 19567 11645 19579 11679
rect 19521 11639 19579 11645
rect 19536 11608 19564 11639
rect 19610 11636 19616 11688
rect 19668 11676 19674 11688
rect 19981 11679 20039 11685
rect 19981 11676 19993 11679
rect 19668 11648 19993 11676
rect 19668 11636 19674 11648
rect 19981 11645 19993 11648
rect 20027 11645 20039 11679
rect 19981 11639 20039 11645
rect 20165 11679 20223 11685
rect 20165 11645 20177 11679
rect 20211 11676 20223 11679
rect 20714 11676 20720 11688
rect 20211 11648 20720 11676
rect 20211 11645 20223 11648
rect 20165 11639 20223 11645
rect 20180 11608 20208 11639
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 19536 11580 20208 11608
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 18325 11543 18383 11549
rect 18325 11540 18337 11543
rect 18104 11512 18337 11540
rect 18104 11500 18110 11512
rect 18325 11509 18337 11512
rect 18371 11509 18383 11543
rect 20438 11540 20444 11552
rect 20399 11512 20444 11540
rect 18325 11503 18383 11509
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 1104 11450 21712 11472
rect 1104 11398 7851 11450
rect 7903 11398 7915 11450
rect 7967 11398 7979 11450
rect 8031 11398 8043 11450
rect 8095 11398 14720 11450
rect 14772 11398 14784 11450
rect 14836 11398 14848 11450
rect 14900 11398 14912 11450
rect 14964 11398 21712 11450
rect 1104 11376 21712 11398
rect 16758 11336 16764 11348
rect 16719 11308 16764 11336
rect 16758 11296 16764 11308
rect 16816 11296 16822 11348
rect 17862 11336 17868 11348
rect 17823 11308 17868 11336
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 18785 11271 18843 11277
rect 18785 11268 18797 11271
rect 13464 11240 18797 11268
rect 13464 11212 13492 11240
rect 18785 11237 18797 11240
rect 18831 11237 18843 11271
rect 18785 11231 18843 11237
rect 10781 11203 10839 11209
rect 10781 11169 10793 11203
rect 10827 11200 10839 11203
rect 11054 11200 11060 11212
rect 10827 11172 11060 11200
rect 10827 11169 10839 11172
rect 10781 11163 10839 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 12345 11203 12403 11209
rect 12345 11169 12357 11203
rect 12391 11200 12403 11203
rect 13446 11200 13452 11212
rect 12391 11172 13452 11200
rect 12391 11169 12403 11172
rect 12345 11163 12403 11169
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 16577 11203 16635 11209
rect 16577 11169 16589 11203
rect 16623 11169 16635 11203
rect 17678 11200 17684 11212
rect 17639 11172 17684 11200
rect 16577 11163 16635 11169
rect 16592 11132 16620 11163
rect 17678 11160 17684 11172
rect 17736 11160 17742 11212
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 19429 11203 19487 11209
rect 19429 11200 19441 11203
rect 19392 11172 19441 11200
rect 19392 11160 19398 11172
rect 19429 11169 19441 11172
rect 19475 11169 19487 11203
rect 19429 11163 19487 11169
rect 19610 11160 19616 11212
rect 19668 11200 19674 11212
rect 19797 11203 19855 11209
rect 19797 11200 19809 11203
rect 19668 11172 19809 11200
rect 19668 11160 19674 11172
rect 19797 11169 19809 11172
rect 19843 11169 19855 11203
rect 19797 11163 19855 11169
rect 19981 11203 20039 11209
rect 19981 11169 19993 11203
rect 20027 11200 20039 11203
rect 20714 11200 20720 11212
rect 20027 11172 20720 11200
rect 20027 11169 20039 11172
rect 19981 11163 20039 11169
rect 20714 11160 20720 11172
rect 20772 11160 20778 11212
rect 19352 11132 19380 11160
rect 19518 11132 19524 11144
rect 16592 11104 19380 11132
rect 19479 11104 19524 11132
rect 19518 11092 19524 11104
rect 19576 11092 19582 11144
rect 10778 11024 10784 11076
rect 10836 11064 10842 11076
rect 10965 11067 11023 11073
rect 10965 11064 10977 11067
rect 10836 11036 10977 11064
rect 10836 11024 10842 11036
rect 10965 11033 10977 11036
rect 11011 11033 11023 11067
rect 10965 11027 11023 11033
rect 12529 10999 12587 11005
rect 12529 10965 12541 10999
rect 12575 10996 12587 10999
rect 12802 10996 12808 11008
rect 12575 10968 12808 10996
rect 12575 10965 12587 10968
rect 12529 10959 12587 10965
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 13633 10999 13691 11005
rect 13633 10996 13645 10999
rect 13412 10968 13645 10996
rect 13412 10956 13418 10968
rect 13633 10965 13645 10968
rect 13679 10965 13691 10999
rect 13633 10959 13691 10965
rect 1104 10906 21712 10928
rect 1104 10854 4416 10906
rect 4468 10854 4480 10906
rect 4532 10854 4544 10906
rect 4596 10854 4608 10906
rect 4660 10854 11286 10906
rect 11338 10854 11350 10906
rect 11402 10854 11414 10906
rect 11466 10854 11478 10906
rect 11530 10854 18155 10906
rect 18207 10854 18219 10906
rect 18271 10854 18283 10906
rect 18335 10854 18347 10906
rect 18399 10854 21712 10906
rect 1104 10832 21712 10854
rect 13817 10795 13875 10801
rect 13817 10761 13829 10795
rect 13863 10792 13875 10795
rect 15194 10792 15200 10804
rect 13863 10764 15200 10792
rect 13863 10761 13875 10764
rect 13817 10755 13875 10761
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 13906 10684 13912 10736
rect 13964 10724 13970 10736
rect 13964 10696 15884 10724
rect 13964 10684 13970 10696
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10656 10563 10659
rect 10594 10656 10600 10668
rect 10551 10628 10600 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 11054 10656 11060 10668
rect 10704 10628 11060 10656
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10588 10471 10591
rect 10704 10588 10732 10628
rect 11054 10616 11060 10628
rect 11112 10656 11118 10668
rect 11790 10656 11796 10668
rect 11112 10628 11796 10656
rect 11112 10616 11118 10628
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 14090 10616 14096 10668
rect 14148 10656 14154 10668
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 14148 10628 15761 10656
rect 14148 10616 14154 10628
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 10459 10560 10732 10588
rect 10781 10591 10839 10597
rect 10459 10557 10471 10560
rect 10413 10551 10471 10557
rect 10781 10557 10793 10591
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 10226 10480 10232 10532
rect 10284 10520 10290 10532
rect 10796 10520 10824 10551
rect 10870 10548 10876 10600
rect 10928 10588 10934 10600
rect 12802 10588 12808 10600
rect 10928 10560 10973 10588
rect 12763 10560 12808 10588
rect 10928 10548 10934 10560
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 12894 10548 12900 10600
rect 12952 10588 12958 10600
rect 13265 10591 13323 10597
rect 13265 10588 13277 10591
rect 12952 10560 13277 10588
rect 12952 10548 12958 10560
rect 13265 10557 13277 10560
rect 13311 10557 13323 10591
rect 13265 10551 13323 10557
rect 13354 10548 13360 10600
rect 13412 10588 13418 10600
rect 13412 10560 13457 10588
rect 13412 10548 13418 10560
rect 14366 10548 14372 10600
rect 14424 10588 14430 10600
rect 15856 10597 15884 10696
rect 19352 10696 20392 10724
rect 19352 10665 19380 10696
rect 19337 10659 19395 10665
rect 19337 10625 19349 10659
rect 19383 10625 19395 10659
rect 19337 10619 19395 10625
rect 15289 10591 15347 10597
rect 15289 10588 15301 10591
rect 14424 10560 15301 10588
rect 14424 10548 14430 10560
rect 15289 10557 15301 10560
rect 15335 10557 15347 10591
rect 15289 10551 15347 10557
rect 15473 10591 15531 10597
rect 15473 10557 15485 10591
rect 15519 10557 15531 10591
rect 15473 10551 15531 10557
rect 15841 10591 15899 10597
rect 15841 10557 15853 10591
rect 15887 10557 15899 10591
rect 15841 10551 15899 10557
rect 15194 10520 15200 10532
rect 10284 10492 10824 10520
rect 15028 10492 15200 10520
rect 10284 10480 10290 10492
rect 10045 10455 10103 10461
rect 10045 10421 10057 10455
rect 10091 10452 10103 10455
rect 15028 10452 15056 10492
rect 15194 10480 15200 10492
rect 15252 10520 15258 10532
rect 15488 10520 15516 10551
rect 18046 10548 18052 10600
rect 18104 10588 18110 10600
rect 18141 10591 18199 10597
rect 18141 10588 18153 10591
rect 18104 10560 18153 10588
rect 18104 10548 18110 10560
rect 18141 10557 18153 10560
rect 18187 10557 18199 10591
rect 19426 10588 19432 10600
rect 19387 10560 19432 10588
rect 18141 10551 18199 10557
rect 19426 10548 19432 10560
rect 19484 10548 19490 10600
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10557 20039 10591
rect 19981 10551 20039 10557
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10588 20223 10591
rect 20364 10588 20392 10696
rect 20438 10588 20444 10600
rect 20211 10560 20444 10588
rect 20211 10557 20223 10560
rect 20165 10551 20223 10557
rect 19996 10520 20024 10551
rect 20438 10548 20444 10560
rect 20496 10548 20502 10600
rect 15252 10492 15516 10520
rect 18340 10492 20024 10520
rect 15252 10480 15258 10492
rect 10091 10424 15056 10452
rect 15105 10455 15163 10461
rect 10091 10421 10103 10424
rect 10045 10415 10103 10421
rect 15105 10421 15117 10455
rect 15151 10452 15163 10455
rect 16574 10452 16580 10464
rect 15151 10424 16580 10452
rect 15151 10421 15163 10424
rect 15105 10415 15163 10421
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 18340 10461 18368 10492
rect 18325 10455 18383 10461
rect 18325 10421 18337 10455
rect 18371 10421 18383 10455
rect 20438 10452 20444 10464
rect 20399 10424 20444 10452
rect 18325 10415 18383 10421
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 1104 10362 21712 10384
rect 1104 10310 7851 10362
rect 7903 10310 7915 10362
rect 7967 10310 7979 10362
rect 8031 10310 8043 10362
rect 8095 10310 14720 10362
rect 14772 10310 14784 10362
rect 14836 10310 14848 10362
rect 14900 10310 14912 10362
rect 14964 10310 21712 10362
rect 1104 10288 21712 10310
rect 19061 10251 19119 10257
rect 19061 10217 19073 10251
rect 19107 10248 19119 10251
rect 19242 10248 19248 10260
rect 19107 10220 19248 10248
rect 19107 10217 19119 10220
rect 19061 10211 19119 10217
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 10594 10180 10600 10192
rect 10555 10152 10600 10180
rect 10594 10140 10600 10152
rect 10652 10140 10658 10192
rect 12805 10183 12863 10189
rect 11532 10152 12388 10180
rect 10137 10115 10195 10121
rect 10137 10081 10149 10115
rect 10183 10112 10195 10115
rect 10226 10112 10232 10124
rect 10183 10084 10232 10112
rect 10183 10081 10195 10084
rect 10137 10075 10195 10081
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 11532 10121 11560 10152
rect 12360 10124 12388 10152
rect 12805 10149 12817 10183
rect 12851 10180 12863 10183
rect 12894 10180 12900 10192
rect 12851 10152 12900 10180
rect 12851 10149 12863 10152
rect 12805 10143 12863 10149
rect 12894 10140 12900 10152
rect 12952 10140 12958 10192
rect 14366 10180 14372 10192
rect 14327 10152 14372 10180
rect 14366 10140 14372 10152
rect 14424 10140 14430 10192
rect 15304 10152 16068 10180
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10081 11575 10115
rect 11517 10075 11575 10081
rect 11606 10072 11612 10124
rect 11664 10112 11670 10124
rect 11701 10115 11759 10121
rect 11701 10112 11713 10115
rect 11664 10084 11713 10112
rect 11664 10072 11670 10084
rect 11701 10081 11713 10084
rect 11747 10112 11759 10115
rect 12253 10115 12311 10121
rect 12253 10112 12265 10115
rect 11747 10084 12265 10112
rect 11747 10081 11759 10084
rect 11701 10075 11759 10081
rect 12253 10081 12265 10084
rect 12299 10081 12311 10115
rect 12253 10075 12311 10081
rect 12342 10072 12348 10124
rect 12400 10112 12406 10124
rect 12437 10115 12495 10121
rect 12437 10112 12449 10115
rect 12400 10084 12449 10112
rect 12400 10072 12406 10084
rect 12437 10081 12449 10084
rect 12483 10081 12495 10115
rect 13906 10112 13912 10124
rect 13867 10084 13912 10112
rect 12437 10075 12495 10081
rect 13906 10072 13912 10084
rect 13964 10072 13970 10124
rect 15194 10072 15200 10124
rect 15252 10112 15258 10124
rect 15304 10121 15332 10152
rect 15289 10115 15347 10121
rect 15289 10112 15301 10115
rect 15252 10084 15301 10112
rect 15252 10072 15258 10084
rect 15289 10081 15301 10084
rect 15335 10081 15347 10115
rect 15470 10112 15476 10124
rect 15431 10084 15476 10112
rect 15289 10075 15347 10081
rect 15470 10072 15476 10084
rect 15528 10112 15534 10124
rect 16040 10121 16068 10152
rect 15933 10115 15991 10121
rect 15933 10112 15945 10115
rect 15528 10084 15945 10112
rect 15528 10072 15534 10084
rect 15933 10081 15945 10084
rect 15979 10081 15991 10115
rect 15933 10075 15991 10081
rect 16025 10115 16083 10121
rect 16025 10081 16037 10115
rect 16071 10081 16083 10115
rect 16025 10075 16083 10081
rect 17586 10072 17592 10124
rect 17644 10112 17650 10124
rect 17681 10115 17739 10121
rect 17681 10112 17693 10115
rect 17644 10084 17693 10112
rect 17644 10072 17650 10084
rect 17681 10081 17693 10084
rect 17727 10112 17739 10115
rect 19429 10115 19487 10121
rect 19429 10112 19441 10115
rect 17727 10084 19441 10112
rect 17727 10081 17739 10084
rect 17681 10075 17739 10081
rect 19429 10081 19441 10084
rect 19475 10081 19487 10115
rect 19429 10075 19487 10081
rect 19797 10115 19855 10121
rect 19797 10081 19809 10115
rect 19843 10112 19855 10115
rect 19978 10112 19984 10124
rect 19843 10084 19984 10112
rect 19843 10081 19855 10084
rect 19797 10075 19855 10081
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 10045 10047 10103 10053
rect 10045 10013 10057 10047
rect 10091 10044 10103 10047
rect 10870 10044 10876 10056
rect 10091 10016 10876 10044
rect 10091 10013 10103 10016
rect 10045 10007 10103 10013
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 13817 10047 13875 10053
rect 13817 10013 13829 10047
rect 13863 10044 13875 10047
rect 14090 10044 14096 10056
rect 13863 10016 14096 10044
rect 13863 10013 13875 10016
rect 13817 10007 13875 10013
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 19518 10044 19524 10056
rect 19479 10016 19524 10044
rect 19518 10004 19524 10016
rect 19576 10004 19582 10056
rect 19702 10044 19708 10056
rect 19663 10016 19708 10044
rect 19702 10004 19708 10016
rect 19760 10004 19766 10056
rect 15102 9936 15108 9988
rect 15160 9976 15166 9988
rect 16393 9979 16451 9985
rect 16393 9976 16405 9979
rect 15160 9948 16405 9976
rect 15160 9936 15166 9948
rect 16393 9945 16405 9948
rect 16439 9945 16451 9979
rect 16393 9939 16451 9945
rect 17865 9911 17923 9917
rect 17865 9877 17877 9911
rect 17911 9908 17923 9911
rect 19058 9908 19064 9920
rect 17911 9880 19064 9908
rect 17911 9877 17923 9880
rect 17865 9871 17923 9877
rect 19058 9868 19064 9880
rect 19116 9868 19122 9920
rect 1104 9818 21712 9840
rect 1104 9766 4416 9818
rect 4468 9766 4480 9818
rect 4532 9766 4544 9818
rect 4596 9766 4608 9818
rect 4660 9766 11286 9818
rect 11338 9766 11350 9818
rect 11402 9766 11414 9818
rect 11466 9766 11478 9818
rect 11530 9766 18155 9818
rect 18207 9766 18219 9818
rect 18271 9766 18283 9818
rect 18335 9766 18347 9818
rect 18399 9766 21712 9818
rect 1104 9744 21712 9766
rect 20162 9636 20168 9648
rect 19628 9608 20168 9636
rect 15105 9571 15163 9577
rect 9876 9540 10088 9568
rect 4062 9460 4068 9512
rect 4120 9500 4126 9512
rect 9876 9509 9904 9540
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 4120 9472 9873 9500
rect 4120 9460 4126 9472
rect 9861 9469 9873 9472
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 9953 9503 10011 9509
rect 9953 9469 9965 9503
rect 9999 9469 10011 9503
rect 10060 9500 10088 9540
rect 15105 9537 15117 9571
rect 15151 9568 15163 9571
rect 15470 9568 15476 9580
rect 15151 9540 15476 9568
rect 15151 9537 15163 9540
rect 15105 9531 15163 9537
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 10226 9500 10232 9512
rect 10060 9472 10232 9500
rect 9953 9463 10011 9469
rect 9968 9432 9996 9463
rect 10226 9460 10232 9472
rect 10284 9500 10290 9512
rect 10413 9503 10471 9509
rect 10413 9500 10425 9503
rect 10284 9472 10425 9500
rect 10284 9460 10290 9472
rect 10413 9469 10425 9472
rect 10459 9469 10471 9503
rect 10413 9463 10471 9469
rect 10597 9503 10655 9509
rect 10597 9469 10609 9503
rect 10643 9500 10655 9503
rect 10870 9500 10876 9512
rect 10643 9472 10876 9500
rect 10643 9469 10655 9472
rect 10597 9463 10655 9469
rect 10612 9432 10640 9463
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 12250 9460 12256 9512
rect 12308 9500 12314 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12308 9472 12449 9500
rect 12308 9460 12314 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 12529 9503 12587 9509
rect 12529 9469 12541 9503
rect 12575 9469 12587 9503
rect 12529 9463 12587 9469
rect 9968 9404 10640 9432
rect 12342 9392 12348 9444
rect 12400 9432 12406 9444
rect 12544 9432 12572 9463
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 14001 9503 14059 9509
rect 14001 9500 14013 9503
rect 13964 9472 14013 9500
rect 13964 9460 13970 9472
rect 14001 9469 14013 9472
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 12400 9404 12572 9432
rect 12989 9435 13047 9441
rect 12400 9392 12406 9404
rect 12989 9401 13001 9435
rect 13035 9432 13047 9435
rect 13262 9432 13268 9444
rect 13035 9404 13268 9432
rect 13035 9401 13047 9404
rect 12989 9395 13047 9401
rect 13262 9392 13268 9404
rect 13320 9392 13326 9444
rect 14016 9432 14044 9463
rect 14090 9460 14096 9512
rect 14148 9500 14154 9512
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14148 9472 14473 9500
rect 14148 9460 14154 9472
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 14553 9503 14611 9509
rect 14553 9469 14565 9503
rect 14599 9469 14611 9503
rect 14553 9463 14611 9469
rect 14568 9432 14596 9463
rect 19058 9460 19064 9512
rect 19116 9500 19122 9512
rect 19429 9503 19487 9509
rect 19429 9500 19441 9503
rect 19116 9472 19441 9500
rect 19116 9460 19122 9472
rect 19429 9469 19441 9472
rect 19475 9469 19487 9503
rect 19429 9463 19487 9469
rect 19521 9503 19579 9509
rect 19521 9469 19533 9503
rect 19567 9500 19579 9503
rect 19628 9500 19656 9608
rect 20162 9596 20168 9608
rect 20220 9596 20226 9648
rect 19979 9503 20037 9509
rect 19979 9500 19991 9503
rect 19567 9472 19656 9500
rect 19720 9472 19991 9500
rect 19567 9469 19579 9472
rect 19521 9463 19579 9469
rect 14016 9404 14596 9432
rect 19444 9432 19472 9463
rect 19720 9432 19748 9472
rect 19979 9469 19991 9472
rect 20025 9469 20037 9503
rect 20162 9500 20168 9512
rect 20123 9472 20168 9500
rect 19979 9463 20037 9469
rect 20162 9460 20168 9472
rect 20220 9460 20226 9512
rect 19444 9404 19748 9432
rect 10870 9364 10876 9376
rect 10831 9336 10876 9364
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 20346 9324 20352 9376
rect 20404 9364 20410 9376
rect 20441 9367 20499 9373
rect 20441 9364 20453 9367
rect 20404 9336 20453 9364
rect 20404 9324 20410 9336
rect 20441 9333 20453 9336
rect 20487 9333 20499 9367
rect 20441 9327 20499 9333
rect 1104 9274 21712 9296
rect 1104 9222 7851 9274
rect 7903 9222 7915 9274
rect 7967 9222 7979 9274
rect 8031 9222 8043 9274
rect 8095 9222 14720 9274
rect 14772 9222 14784 9274
rect 14836 9222 14848 9274
rect 14900 9222 14912 9274
rect 14964 9222 21712 9274
rect 1104 9200 21712 9222
rect 10888 9064 11560 9092
rect 10888 9036 10916 9064
rect 10778 9024 10784 9036
rect 10739 8996 10784 9024
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 10928 8996 10973 9024
rect 10928 8984 10934 8996
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 11532 9033 11560 9064
rect 11606 9052 11612 9104
rect 11664 9092 11670 9104
rect 12342 9092 12348 9104
rect 11664 9064 12348 9092
rect 11664 9052 11670 9064
rect 12342 9052 12348 9064
rect 12400 9092 12406 9104
rect 12400 9064 13860 9092
rect 12400 9052 12406 9064
rect 11333 9027 11391 9033
rect 11333 9024 11345 9027
rect 11204 8996 11345 9024
rect 11204 8984 11210 8996
rect 11333 8993 11345 8996
rect 11379 8993 11391 9027
rect 11333 8987 11391 8993
rect 11517 9027 11575 9033
rect 11517 8993 11529 9027
rect 11563 8993 11575 9027
rect 13262 9024 13268 9036
rect 13223 8996 13268 9024
rect 11517 8987 11575 8993
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 13446 9024 13452 9036
rect 13407 8996 13452 9024
rect 13446 8984 13452 8996
rect 13504 8984 13510 9036
rect 13832 9033 13860 9064
rect 13817 9027 13875 9033
rect 13817 8993 13829 9027
rect 13863 8993 13875 9027
rect 13817 8987 13875 8993
rect 19521 9027 19579 9033
rect 19521 8993 19533 9027
rect 19567 9024 19579 9027
rect 19978 9024 19984 9036
rect 19567 8996 19984 9024
rect 19567 8993 19579 8996
rect 19521 8987 19579 8993
rect 19978 8984 19984 8996
rect 20036 8984 20042 9036
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 11848 8928 12817 8956
rect 11848 8916 11854 8928
rect 12805 8925 12817 8928
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8956 19487 8959
rect 19702 8956 19708 8968
rect 19475 8928 19708 8956
rect 19475 8925 19487 8928
rect 19429 8919 19487 8925
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 12250 8888 12256 8900
rect 11756 8860 12256 8888
rect 11756 8848 11762 8860
rect 12250 8848 12256 8860
rect 12308 8888 12314 8900
rect 13740 8888 13768 8919
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 12308 8860 13768 8888
rect 12308 8848 12314 8860
rect 11793 8823 11851 8829
rect 11793 8789 11805 8823
rect 11839 8820 11851 8823
rect 11974 8820 11980 8832
rect 11839 8792 11980 8820
rect 11839 8789 11851 8792
rect 11793 8783 11851 8789
rect 11974 8780 11980 8792
rect 12032 8780 12038 8832
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 19705 8823 19763 8829
rect 19705 8820 19717 8823
rect 19576 8792 19717 8820
rect 19576 8780 19582 8792
rect 19705 8789 19717 8792
rect 19751 8789 19763 8823
rect 19705 8783 19763 8789
rect 1104 8730 21712 8752
rect 1104 8678 4416 8730
rect 4468 8678 4480 8730
rect 4532 8678 4544 8730
rect 4596 8678 4608 8730
rect 4660 8678 11286 8730
rect 11338 8678 11350 8730
rect 11402 8678 11414 8730
rect 11466 8678 11478 8730
rect 11530 8678 18155 8730
rect 18207 8678 18219 8730
rect 18271 8678 18283 8730
rect 18335 8678 18347 8730
rect 18399 8678 21712 8730
rect 1104 8656 21712 8678
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 11425 8619 11483 8625
rect 11425 8616 11437 8619
rect 11204 8588 11437 8616
rect 11204 8576 11210 8588
rect 11425 8585 11437 8588
rect 11471 8585 11483 8619
rect 11425 8579 11483 8585
rect 20162 8508 20168 8560
rect 20220 8548 20226 8560
rect 20349 8551 20407 8557
rect 20349 8548 20361 8551
rect 20220 8520 20361 8548
rect 20220 8508 20226 8520
rect 20349 8517 20361 8520
rect 20395 8517 20407 8551
rect 20349 8511 20407 8517
rect 11241 8415 11299 8421
rect 11241 8381 11253 8415
rect 11287 8412 11299 8415
rect 11790 8412 11796 8424
rect 11287 8384 11796 8412
rect 11287 8381 11299 8384
rect 11241 8375 11299 8381
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 19429 8415 19487 8421
rect 19429 8381 19441 8415
rect 19475 8381 19487 8415
rect 19429 8375 19487 8381
rect 19521 8415 19579 8421
rect 19521 8381 19533 8415
rect 19567 8412 19579 8415
rect 19610 8412 19616 8424
rect 19567 8384 19616 8412
rect 19567 8381 19579 8384
rect 19521 8375 19579 8381
rect 19444 8344 19472 8375
rect 19610 8372 19616 8384
rect 19668 8412 19674 8424
rect 19889 8415 19947 8421
rect 19889 8412 19901 8415
rect 19668 8384 19901 8412
rect 19668 8372 19674 8384
rect 19889 8381 19901 8384
rect 19935 8381 19947 8415
rect 19889 8375 19947 8381
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 20036 8384 20081 8412
rect 20036 8372 20042 8384
rect 19996 8344 20024 8372
rect 19444 8316 20024 8344
rect 1104 8186 21712 8208
rect 1104 8134 7851 8186
rect 7903 8134 7915 8186
rect 7967 8134 7979 8186
rect 8031 8134 8043 8186
rect 8095 8134 14720 8186
rect 14772 8134 14784 8186
rect 14836 8134 14848 8186
rect 14900 8134 14912 8186
rect 14964 8134 21712 8186
rect 1104 8112 21712 8134
rect 1104 7642 21712 7664
rect 1104 7590 4416 7642
rect 4468 7590 4480 7642
rect 4532 7590 4544 7642
rect 4596 7590 4608 7642
rect 4660 7590 11286 7642
rect 11338 7590 11350 7642
rect 11402 7590 11414 7642
rect 11466 7590 11478 7642
rect 11530 7590 18155 7642
rect 18207 7590 18219 7642
rect 18271 7590 18283 7642
rect 18335 7590 18347 7642
rect 18399 7590 21712 7642
rect 1104 7568 21712 7590
rect 1104 7098 21712 7120
rect 1104 7046 7851 7098
rect 7903 7046 7915 7098
rect 7967 7046 7979 7098
rect 8031 7046 8043 7098
rect 8095 7046 14720 7098
rect 14772 7046 14784 7098
rect 14836 7046 14848 7098
rect 14900 7046 14912 7098
rect 14964 7046 21712 7098
rect 1104 7024 21712 7046
rect 1104 6554 21712 6576
rect 1104 6502 4416 6554
rect 4468 6502 4480 6554
rect 4532 6502 4544 6554
rect 4596 6502 4608 6554
rect 4660 6502 11286 6554
rect 11338 6502 11350 6554
rect 11402 6502 11414 6554
rect 11466 6502 11478 6554
rect 11530 6502 18155 6554
rect 18207 6502 18219 6554
rect 18271 6502 18283 6554
rect 18335 6502 18347 6554
rect 18399 6502 21712 6554
rect 1104 6480 21712 6502
rect 1104 6010 21712 6032
rect 1104 5958 7851 6010
rect 7903 5958 7915 6010
rect 7967 5958 7979 6010
rect 8031 5958 8043 6010
rect 8095 5958 14720 6010
rect 14772 5958 14784 6010
rect 14836 5958 14848 6010
rect 14900 5958 14912 6010
rect 14964 5958 21712 6010
rect 1104 5936 21712 5958
rect 1104 5466 21712 5488
rect 1104 5414 4416 5466
rect 4468 5414 4480 5466
rect 4532 5414 4544 5466
rect 4596 5414 4608 5466
rect 4660 5414 11286 5466
rect 11338 5414 11350 5466
rect 11402 5414 11414 5466
rect 11466 5414 11478 5466
rect 11530 5414 18155 5466
rect 18207 5414 18219 5466
rect 18271 5414 18283 5466
rect 18335 5414 18347 5466
rect 18399 5414 21712 5466
rect 1104 5392 21712 5414
rect 1104 4922 21712 4944
rect 1104 4870 7851 4922
rect 7903 4870 7915 4922
rect 7967 4870 7979 4922
rect 8031 4870 8043 4922
rect 8095 4870 14720 4922
rect 14772 4870 14784 4922
rect 14836 4870 14848 4922
rect 14900 4870 14912 4922
rect 14964 4870 21712 4922
rect 1104 4848 21712 4870
rect 1104 4378 21712 4400
rect 1104 4326 4416 4378
rect 4468 4326 4480 4378
rect 4532 4326 4544 4378
rect 4596 4326 4608 4378
rect 4660 4326 11286 4378
rect 11338 4326 11350 4378
rect 11402 4326 11414 4378
rect 11466 4326 11478 4378
rect 11530 4326 18155 4378
rect 18207 4326 18219 4378
rect 18271 4326 18283 4378
rect 18335 4326 18347 4378
rect 18399 4326 21712 4378
rect 1104 4304 21712 4326
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 11606 4128 11612 4140
rect 9272 4100 11612 4128
rect 9272 4088 9278 4100
rect 11606 4088 11612 4100
rect 11664 4088 11670 4140
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 11698 4060 11704 4072
rect 6328 4032 11704 4060
rect 6328 4020 6334 4032
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 1104 3834 21712 3856
rect 1104 3782 7851 3834
rect 7903 3782 7915 3834
rect 7967 3782 7979 3834
rect 8031 3782 8043 3834
rect 8095 3782 14720 3834
rect 14772 3782 14784 3834
rect 14836 3782 14848 3834
rect 14900 3782 14912 3834
rect 14964 3782 21712 3834
rect 1104 3760 21712 3782
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1486 3516 1492 3528
rect 624 3488 1492 3516
rect 624 3476 630 3488
rect 1486 3476 1492 3488
rect 1544 3476 1550 3528
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 17862 3516 17868 3528
rect 16632 3488 17868 3516
rect 16632 3476 16638 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 1104 3290 21712 3312
rect 1104 3238 4416 3290
rect 4468 3238 4480 3290
rect 4532 3238 4544 3290
rect 4596 3238 4608 3290
rect 4660 3238 11286 3290
rect 11338 3238 11350 3290
rect 11402 3238 11414 3290
rect 11466 3238 11478 3290
rect 11530 3238 18155 3290
rect 18207 3238 18219 3290
rect 18271 3238 18283 3290
rect 18335 3238 18347 3290
rect 18399 3238 21712 3290
rect 1104 3216 21712 3238
rect 1104 2746 21712 2768
rect 1104 2694 7851 2746
rect 7903 2694 7915 2746
rect 7967 2694 7979 2746
rect 8031 2694 8043 2746
rect 8095 2694 14720 2746
rect 14772 2694 14784 2746
rect 14836 2694 14848 2746
rect 14900 2694 14912 2746
rect 14964 2694 21712 2746
rect 1104 2672 21712 2694
rect 1104 2202 21712 2224
rect 1104 2150 4416 2202
rect 4468 2150 4480 2202
rect 4532 2150 4544 2202
rect 4596 2150 4608 2202
rect 4660 2150 11286 2202
rect 11338 2150 11350 2202
rect 11402 2150 11414 2202
rect 11466 2150 11478 2202
rect 11530 2150 18155 2202
rect 18207 2150 18219 2202
rect 18271 2150 18283 2202
rect 18335 2150 18347 2202
rect 18399 2150 21712 2202
rect 1104 2128 21712 2150
<< via1 >>
rect 7851 22278 7903 22330
rect 7915 22278 7967 22330
rect 7979 22278 8031 22330
rect 8043 22278 8095 22330
rect 14720 22278 14772 22330
rect 14784 22278 14836 22330
rect 14848 22278 14900 22330
rect 14912 22278 14964 22330
rect 4252 22040 4304 22092
rect 13176 22040 13228 22092
rect 14556 21972 14608 22024
rect 4712 21836 4764 21888
rect 12992 21879 13044 21888
rect 12992 21845 13001 21879
rect 13001 21845 13035 21879
rect 13035 21845 13044 21879
rect 12992 21836 13044 21845
rect 13820 21836 13872 21888
rect 4416 21734 4468 21786
rect 4480 21734 4532 21786
rect 4544 21734 4596 21786
rect 4608 21734 4660 21786
rect 11286 21734 11338 21786
rect 11350 21734 11402 21786
rect 11414 21734 11466 21786
rect 11478 21734 11530 21786
rect 18155 21734 18207 21786
rect 18219 21734 18271 21786
rect 18283 21734 18335 21786
rect 18347 21734 18399 21786
rect 4804 21632 4856 21684
rect 13452 21632 13504 21684
rect 3148 21471 3200 21480
rect 3148 21437 3157 21471
rect 3157 21437 3191 21471
rect 3191 21437 3200 21471
rect 3148 21428 3200 21437
rect 3332 21471 3384 21480
rect 3332 21437 3341 21471
rect 3341 21437 3375 21471
rect 3375 21437 3384 21471
rect 3332 21428 3384 21437
rect 2044 21292 2096 21344
rect 13084 21471 13136 21480
rect 13084 21437 13093 21471
rect 13093 21437 13127 21471
rect 13127 21437 13136 21471
rect 13084 21428 13136 21437
rect 12992 21360 13044 21412
rect 14096 21360 14148 21412
rect 19340 21360 19392 21412
rect 4068 21292 4120 21344
rect 7851 21190 7903 21242
rect 7915 21190 7967 21242
rect 7979 21190 8031 21242
rect 8043 21190 8095 21242
rect 14720 21190 14772 21242
rect 14784 21190 14836 21242
rect 14848 21190 14900 21242
rect 14912 21190 14964 21242
rect 2228 21088 2280 21140
rect 1584 21020 1636 21072
rect 3332 21088 3384 21140
rect 13084 21088 13136 21140
rect 2044 20995 2096 21004
rect 2044 20961 2053 20995
rect 2053 20961 2087 20995
rect 2087 20961 2096 20995
rect 2044 20952 2096 20961
rect 4068 20995 4120 21004
rect 4068 20961 4077 20995
rect 4077 20961 4111 20995
rect 4111 20961 4120 20995
rect 4068 20952 4120 20961
rect 11888 20952 11940 21004
rect 2136 20927 2188 20936
rect 2136 20893 2145 20927
rect 2145 20893 2179 20927
rect 2179 20893 2188 20927
rect 2136 20884 2188 20893
rect 2320 20927 2372 20936
rect 2320 20893 2329 20927
rect 2329 20893 2363 20927
rect 2363 20893 2372 20927
rect 2320 20884 2372 20893
rect 7748 20884 7800 20936
rect 12440 21020 12492 21072
rect 12716 20995 12768 21004
rect 12716 20961 12725 20995
rect 12725 20961 12759 20995
rect 12759 20961 12768 20995
rect 12716 20952 12768 20961
rect 13360 20952 13412 21004
rect 15292 20995 15344 21004
rect 15292 20961 15301 20995
rect 15301 20961 15335 20995
rect 15335 20961 15344 20995
rect 15292 20952 15344 20961
rect 13084 20816 13136 20868
rect 4252 20791 4304 20800
rect 4252 20757 4261 20791
rect 4261 20757 4295 20791
rect 4295 20757 4304 20791
rect 4252 20748 4304 20757
rect 12808 20748 12860 20800
rect 15476 20791 15528 20800
rect 15476 20757 15485 20791
rect 15485 20757 15519 20791
rect 15519 20757 15528 20791
rect 15476 20748 15528 20757
rect 4416 20646 4468 20698
rect 4480 20646 4532 20698
rect 4544 20646 4596 20698
rect 4608 20646 4660 20698
rect 11286 20646 11338 20698
rect 11350 20646 11402 20698
rect 11414 20646 11466 20698
rect 11478 20646 11530 20698
rect 18155 20646 18207 20698
rect 18219 20646 18271 20698
rect 18283 20646 18335 20698
rect 18347 20646 18399 20698
rect 12716 20544 12768 20596
rect 1492 20451 1544 20460
rect 1492 20417 1501 20451
rect 1501 20417 1535 20451
rect 1535 20417 1544 20451
rect 2320 20476 2372 20528
rect 4252 20476 4304 20528
rect 14556 20544 14608 20596
rect 12992 20451 13044 20460
rect 1492 20408 1544 20417
rect 1584 20383 1636 20392
rect 1584 20349 1593 20383
rect 1593 20349 1627 20383
rect 1627 20349 1636 20383
rect 1584 20340 1636 20349
rect 12992 20417 13001 20451
rect 13001 20417 13035 20451
rect 13035 20417 13044 20451
rect 12992 20408 13044 20417
rect 13360 20451 13412 20460
rect 13360 20417 13369 20451
rect 13369 20417 13403 20451
rect 13403 20417 13412 20451
rect 13360 20408 13412 20417
rect 3608 20383 3660 20392
rect 3608 20349 3617 20383
rect 3617 20349 3651 20383
rect 3651 20349 3660 20383
rect 3608 20340 3660 20349
rect 4712 20383 4764 20392
rect 4712 20349 4721 20383
rect 4721 20349 4755 20383
rect 4755 20349 4764 20383
rect 4712 20340 4764 20349
rect 13084 20383 13136 20392
rect 13084 20349 13093 20383
rect 13093 20349 13127 20383
rect 13127 20349 13136 20383
rect 13084 20340 13136 20349
rect 15200 20408 15252 20460
rect 16396 20408 16448 20460
rect 18420 20408 18472 20460
rect 20720 20408 20772 20460
rect 22100 20408 22152 20460
rect 15476 20340 15528 20392
rect 2596 20247 2648 20256
rect 2596 20213 2605 20247
rect 2605 20213 2639 20247
rect 2639 20213 2648 20247
rect 2596 20204 2648 20213
rect 4068 20204 4120 20256
rect 17684 20204 17736 20256
rect 7851 20102 7903 20154
rect 7915 20102 7967 20154
rect 7979 20102 8031 20154
rect 8043 20102 8095 20154
rect 14720 20102 14772 20154
rect 14784 20102 14836 20154
rect 14848 20102 14900 20154
rect 14912 20102 14964 20154
rect 3608 20000 3660 20052
rect 11888 20000 11940 20052
rect 2136 19932 2188 19984
rect 12992 19975 13044 19984
rect 12992 19941 13001 19975
rect 13001 19941 13035 19975
rect 13035 19941 13044 19975
rect 12992 19932 13044 19941
rect 1584 19864 1636 19916
rect 4068 19907 4120 19916
rect 4068 19873 4077 19907
rect 4077 19873 4111 19907
rect 4111 19873 4120 19907
rect 4068 19864 4120 19873
rect 12440 19907 12492 19916
rect 12440 19873 12449 19907
rect 12449 19873 12483 19907
rect 12483 19873 12492 19907
rect 12440 19864 12492 19873
rect 12716 19864 12768 19916
rect 13820 19907 13872 19916
rect 13820 19873 13829 19907
rect 13829 19873 13863 19907
rect 13863 19873 13872 19907
rect 13820 19864 13872 19873
rect 1492 19796 1544 19848
rect 4416 19558 4468 19610
rect 4480 19558 4532 19610
rect 4544 19558 4596 19610
rect 4608 19558 4660 19610
rect 11286 19558 11338 19610
rect 11350 19558 11402 19610
rect 11414 19558 11466 19610
rect 11478 19558 11530 19610
rect 18155 19558 18207 19610
rect 18219 19558 18271 19610
rect 18283 19558 18335 19610
rect 18347 19558 18399 19610
rect 4252 19295 4304 19304
rect 4252 19261 4261 19295
rect 4261 19261 4295 19295
rect 4295 19261 4304 19295
rect 4252 19252 4304 19261
rect 6460 19252 6512 19304
rect 12808 19295 12860 19304
rect 12808 19261 12817 19295
rect 12817 19261 12851 19295
rect 12851 19261 12860 19295
rect 12808 19252 12860 19261
rect 1768 19116 1820 19168
rect 2320 19116 2372 19168
rect 4712 19116 4764 19168
rect 15292 19116 15344 19168
rect 7851 19014 7903 19066
rect 7915 19014 7967 19066
rect 7979 19014 8031 19066
rect 8043 19014 8095 19066
rect 14720 19014 14772 19066
rect 14784 19014 14836 19066
rect 14848 19014 14900 19066
rect 14912 19014 14964 19066
rect 6460 18955 6512 18964
rect 6460 18921 6469 18955
rect 6469 18921 6503 18955
rect 6503 18921 6512 18955
rect 6460 18912 6512 18921
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 2320 18776 2372 18828
rect 2596 18776 2648 18828
rect 5172 18819 5224 18828
rect 5172 18785 5181 18819
rect 5181 18785 5215 18819
rect 5215 18785 5224 18819
rect 5172 18776 5224 18785
rect 5264 18776 5316 18828
rect 2688 18615 2740 18624
rect 2688 18581 2697 18615
rect 2697 18581 2731 18615
rect 2731 18581 2740 18615
rect 2688 18572 2740 18581
rect 4252 18615 4304 18624
rect 4252 18581 4261 18615
rect 4261 18581 4295 18615
rect 4295 18581 4304 18615
rect 4252 18572 4304 18581
rect 4416 18470 4468 18522
rect 4480 18470 4532 18522
rect 4544 18470 4596 18522
rect 4608 18470 4660 18522
rect 11286 18470 11338 18522
rect 11350 18470 11402 18522
rect 11414 18470 11466 18522
rect 11478 18470 11530 18522
rect 18155 18470 18207 18522
rect 18219 18470 18271 18522
rect 18283 18470 18335 18522
rect 18347 18470 18399 18522
rect 2044 18368 2096 18420
rect 2228 18232 2280 18284
rect 2504 18207 2556 18216
rect 2504 18173 2513 18207
rect 2513 18173 2547 18207
rect 2547 18173 2556 18207
rect 2504 18164 2556 18173
rect 2780 18164 2832 18216
rect 3056 18207 3108 18216
rect 3056 18173 3065 18207
rect 3065 18173 3099 18207
rect 3099 18173 3108 18207
rect 3056 18164 3108 18173
rect 3148 18164 3200 18216
rect 4160 18164 4212 18216
rect 7851 17926 7903 17978
rect 7915 17926 7967 17978
rect 7979 17926 8031 17978
rect 8043 17926 8095 17978
rect 14720 17926 14772 17978
rect 14784 17926 14836 17978
rect 14848 17926 14900 17978
rect 14912 17926 14964 17978
rect 2504 17756 2556 17808
rect 2780 17688 2832 17740
rect 4712 17688 4764 17740
rect 2872 17620 2924 17672
rect 3056 17620 3108 17672
rect 1584 17527 1636 17536
rect 1584 17493 1593 17527
rect 1593 17493 1627 17527
rect 1627 17493 1636 17527
rect 1584 17484 1636 17493
rect 2504 17484 2556 17536
rect 2872 17484 2924 17536
rect 4416 17382 4468 17434
rect 4480 17382 4532 17434
rect 4544 17382 4596 17434
rect 4608 17382 4660 17434
rect 11286 17382 11338 17434
rect 11350 17382 11402 17434
rect 11414 17382 11466 17434
rect 11478 17382 11530 17434
rect 18155 17382 18207 17434
rect 18219 17382 18271 17434
rect 18283 17382 18335 17434
rect 18347 17382 18399 17434
rect 5172 17280 5224 17332
rect 4160 17212 4212 17264
rect 1584 17144 1636 17196
rect 2872 17076 2924 17128
rect 4252 17008 4304 17060
rect 3976 16983 4028 16992
rect 3976 16949 3985 16983
rect 3985 16949 4019 16983
rect 4019 16949 4028 16983
rect 3976 16940 4028 16949
rect 7851 16838 7903 16890
rect 7915 16838 7967 16890
rect 7979 16838 8031 16890
rect 8043 16838 8095 16890
rect 14720 16838 14772 16890
rect 14784 16838 14836 16890
rect 14848 16838 14900 16890
rect 14912 16838 14964 16890
rect 5264 16736 5316 16788
rect 3976 16600 4028 16652
rect 4416 16294 4468 16346
rect 4480 16294 4532 16346
rect 4544 16294 4596 16346
rect 4608 16294 4660 16346
rect 11286 16294 11338 16346
rect 11350 16294 11402 16346
rect 11414 16294 11466 16346
rect 11478 16294 11530 16346
rect 18155 16294 18207 16346
rect 18219 16294 18271 16346
rect 18283 16294 18335 16346
rect 18347 16294 18399 16346
rect 7851 15750 7903 15802
rect 7915 15750 7967 15802
rect 7979 15750 8031 15802
rect 8043 15750 8095 15802
rect 14720 15750 14772 15802
rect 14784 15750 14836 15802
rect 14848 15750 14900 15802
rect 14912 15750 14964 15802
rect 4416 15206 4468 15258
rect 4480 15206 4532 15258
rect 4544 15206 4596 15258
rect 4608 15206 4660 15258
rect 11286 15206 11338 15258
rect 11350 15206 11402 15258
rect 11414 15206 11466 15258
rect 11478 15206 11530 15258
rect 18155 15206 18207 15258
rect 18219 15206 18271 15258
rect 18283 15206 18335 15258
rect 18347 15206 18399 15258
rect 7851 14662 7903 14714
rect 7915 14662 7967 14714
rect 7979 14662 8031 14714
rect 8043 14662 8095 14714
rect 14720 14662 14772 14714
rect 14784 14662 14836 14714
rect 14848 14662 14900 14714
rect 14912 14662 14964 14714
rect 4416 14118 4468 14170
rect 4480 14118 4532 14170
rect 4544 14118 4596 14170
rect 4608 14118 4660 14170
rect 11286 14118 11338 14170
rect 11350 14118 11402 14170
rect 11414 14118 11466 14170
rect 11478 14118 11530 14170
rect 18155 14118 18207 14170
rect 18219 14118 18271 14170
rect 18283 14118 18335 14170
rect 18347 14118 18399 14170
rect 7851 13574 7903 13626
rect 7915 13574 7967 13626
rect 7979 13574 8031 13626
rect 8043 13574 8095 13626
rect 14720 13574 14772 13626
rect 14784 13574 14836 13626
rect 14848 13574 14900 13626
rect 14912 13574 14964 13626
rect 4416 13030 4468 13082
rect 4480 13030 4532 13082
rect 4544 13030 4596 13082
rect 4608 13030 4660 13082
rect 11286 13030 11338 13082
rect 11350 13030 11402 13082
rect 11414 13030 11466 13082
rect 11478 13030 11530 13082
rect 18155 13030 18207 13082
rect 18219 13030 18271 13082
rect 18283 13030 18335 13082
rect 18347 13030 18399 13082
rect 19340 12724 19392 12776
rect 3424 12588 3476 12640
rect 13912 12588 13964 12640
rect 19432 12588 19484 12640
rect 7851 12486 7903 12538
rect 7915 12486 7967 12538
rect 7979 12486 8031 12538
rect 8043 12486 8095 12538
rect 14720 12486 14772 12538
rect 14784 12486 14836 12538
rect 14848 12486 14900 12538
rect 14912 12486 14964 12538
rect 16764 12248 16816 12300
rect 19524 12291 19576 12300
rect 19524 12257 19533 12291
rect 19533 12257 19567 12291
rect 19567 12257 19576 12291
rect 19524 12248 19576 12257
rect 20720 12180 20772 12232
rect 17684 12044 17736 12096
rect 19524 12044 19576 12096
rect 4416 11942 4468 11994
rect 4480 11942 4532 11994
rect 4544 11942 4596 11994
rect 4608 11942 4660 11994
rect 11286 11942 11338 11994
rect 11350 11942 11402 11994
rect 11414 11942 11466 11994
rect 11478 11942 11530 11994
rect 18155 11942 18207 11994
rect 18219 11942 18271 11994
rect 18283 11942 18335 11994
rect 18347 11942 18399 11994
rect 17868 11636 17920 11688
rect 19616 11636 19668 11688
rect 20720 11636 20772 11688
rect 18052 11500 18104 11552
rect 20444 11543 20496 11552
rect 20444 11509 20453 11543
rect 20453 11509 20487 11543
rect 20487 11509 20496 11543
rect 20444 11500 20496 11509
rect 7851 11398 7903 11450
rect 7915 11398 7967 11450
rect 7979 11398 8031 11450
rect 8043 11398 8095 11450
rect 14720 11398 14772 11450
rect 14784 11398 14836 11450
rect 14848 11398 14900 11450
rect 14912 11398 14964 11450
rect 16764 11339 16816 11348
rect 16764 11305 16773 11339
rect 16773 11305 16807 11339
rect 16807 11305 16816 11339
rect 16764 11296 16816 11305
rect 17868 11339 17920 11348
rect 17868 11305 17877 11339
rect 17877 11305 17911 11339
rect 17911 11305 17920 11339
rect 17868 11296 17920 11305
rect 11060 11160 11112 11212
rect 13452 11203 13504 11212
rect 13452 11169 13461 11203
rect 13461 11169 13495 11203
rect 13495 11169 13504 11203
rect 13452 11160 13504 11169
rect 17684 11203 17736 11212
rect 17684 11169 17693 11203
rect 17693 11169 17727 11203
rect 17727 11169 17736 11203
rect 17684 11160 17736 11169
rect 19340 11160 19392 11212
rect 19616 11160 19668 11212
rect 20720 11160 20772 11212
rect 19524 11135 19576 11144
rect 19524 11101 19533 11135
rect 19533 11101 19567 11135
rect 19567 11101 19576 11135
rect 19524 11092 19576 11101
rect 10784 11024 10836 11076
rect 12808 10956 12860 11008
rect 13360 10956 13412 11008
rect 4416 10854 4468 10906
rect 4480 10854 4532 10906
rect 4544 10854 4596 10906
rect 4608 10854 4660 10906
rect 11286 10854 11338 10906
rect 11350 10854 11402 10906
rect 11414 10854 11466 10906
rect 11478 10854 11530 10906
rect 18155 10854 18207 10906
rect 18219 10854 18271 10906
rect 18283 10854 18335 10906
rect 18347 10854 18399 10906
rect 15200 10752 15252 10804
rect 13912 10684 13964 10736
rect 10600 10616 10652 10668
rect 11060 10616 11112 10668
rect 11796 10616 11848 10668
rect 14096 10616 14148 10668
rect 10232 10480 10284 10532
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 12808 10591 12860 10600
rect 10876 10548 10928 10557
rect 12808 10557 12817 10591
rect 12817 10557 12851 10591
rect 12851 10557 12860 10591
rect 12808 10548 12860 10557
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 13360 10591 13412 10600
rect 13360 10557 13369 10591
rect 13369 10557 13403 10591
rect 13403 10557 13412 10591
rect 13360 10548 13412 10557
rect 14372 10548 14424 10600
rect 15200 10480 15252 10532
rect 18052 10548 18104 10600
rect 19432 10591 19484 10600
rect 19432 10557 19441 10591
rect 19441 10557 19475 10591
rect 19475 10557 19484 10591
rect 19432 10548 19484 10557
rect 20444 10548 20496 10600
rect 16580 10412 16632 10464
rect 20444 10455 20496 10464
rect 20444 10421 20453 10455
rect 20453 10421 20487 10455
rect 20487 10421 20496 10455
rect 20444 10412 20496 10421
rect 7851 10310 7903 10362
rect 7915 10310 7967 10362
rect 7979 10310 8031 10362
rect 8043 10310 8095 10362
rect 14720 10310 14772 10362
rect 14784 10310 14836 10362
rect 14848 10310 14900 10362
rect 14912 10310 14964 10362
rect 19248 10208 19300 10260
rect 10600 10183 10652 10192
rect 10600 10149 10609 10183
rect 10609 10149 10643 10183
rect 10643 10149 10652 10183
rect 10600 10140 10652 10149
rect 10232 10072 10284 10124
rect 12900 10140 12952 10192
rect 14372 10183 14424 10192
rect 14372 10149 14381 10183
rect 14381 10149 14415 10183
rect 14415 10149 14424 10183
rect 14372 10140 14424 10149
rect 11612 10072 11664 10124
rect 12348 10072 12400 10124
rect 13912 10115 13964 10124
rect 13912 10081 13921 10115
rect 13921 10081 13955 10115
rect 13955 10081 13964 10115
rect 13912 10072 13964 10081
rect 15200 10072 15252 10124
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 17592 10072 17644 10124
rect 19984 10072 20036 10124
rect 10876 10004 10928 10056
rect 14096 10004 14148 10056
rect 19524 10047 19576 10056
rect 19524 10013 19533 10047
rect 19533 10013 19567 10047
rect 19567 10013 19576 10047
rect 19524 10004 19576 10013
rect 19708 10047 19760 10056
rect 19708 10013 19717 10047
rect 19717 10013 19751 10047
rect 19751 10013 19760 10047
rect 19708 10004 19760 10013
rect 15108 9936 15160 9988
rect 19064 9868 19116 9920
rect 4416 9766 4468 9818
rect 4480 9766 4532 9818
rect 4544 9766 4596 9818
rect 4608 9766 4660 9818
rect 11286 9766 11338 9818
rect 11350 9766 11402 9818
rect 11414 9766 11466 9818
rect 11478 9766 11530 9818
rect 18155 9766 18207 9818
rect 18219 9766 18271 9818
rect 18283 9766 18335 9818
rect 18347 9766 18399 9818
rect 4068 9460 4120 9512
rect 15476 9528 15528 9580
rect 10232 9460 10284 9512
rect 10876 9460 10928 9512
rect 12256 9460 12308 9512
rect 12348 9392 12400 9444
rect 13912 9460 13964 9512
rect 13268 9392 13320 9444
rect 14096 9503 14148 9512
rect 14096 9469 14105 9503
rect 14105 9469 14139 9503
rect 14139 9469 14148 9503
rect 14096 9460 14148 9469
rect 19064 9460 19116 9512
rect 20168 9596 20220 9648
rect 20168 9503 20220 9512
rect 20168 9469 20177 9503
rect 20177 9469 20211 9503
rect 20211 9469 20220 9503
rect 20168 9460 20220 9469
rect 10876 9367 10928 9376
rect 10876 9333 10885 9367
rect 10885 9333 10919 9367
rect 10919 9333 10928 9367
rect 10876 9324 10928 9333
rect 20352 9324 20404 9376
rect 7851 9222 7903 9274
rect 7915 9222 7967 9274
rect 7979 9222 8031 9274
rect 8043 9222 8095 9274
rect 14720 9222 14772 9274
rect 14784 9222 14836 9274
rect 14848 9222 14900 9274
rect 14912 9222 14964 9274
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 10876 9027 10928 9036
rect 10876 8993 10885 9027
rect 10885 8993 10919 9027
rect 10919 8993 10928 9027
rect 10876 8984 10928 8993
rect 11152 8984 11204 9036
rect 11612 9052 11664 9104
rect 12348 9052 12400 9104
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 13452 9027 13504 9036
rect 13452 8993 13461 9027
rect 13461 8993 13495 9027
rect 13495 8993 13504 9027
rect 13452 8984 13504 8993
rect 19984 8984 20036 9036
rect 11796 8916 11848 8968
rect 11704 8848 11756 8900
rect 12256 8848 12308 8900
rect 19708 8916 19760 8968
rect 11980 8780 12032 8832
rect 19524 8780 19576 8832
rect 4416 8678 4468 8730
rect 4480 8678 4532 8730
rect 4544 8678 4596 8730
rect 4608 8678 4660 8730
rect 11286 8678 11338 8730
rect 11350 8678 11402 8730
rect 11414 8678 11466 8730
rect 11478 8678 11530 8730
rect 18155 8678 18207 8730
rect 18219 8678 18271 8730
rect 18283 8678 18335 8730
rect 18347 8678 18399 8730
rect 11152 8576 11204 8628
rect 20168 8508 20220 8560
rect 11796 8372 11848 8424
rect 19616 8372 19668 8424
rect 19984 8415 20036 8424
rect 19984 8381 19993 8415
rect 19993 8381 20027 8415
rect 20027 8381 20036 8415
rect 19984 8372 20036 8381
rect 7851 8134 7903 8186
rect 7915 8134 7967 8186
rect 7979 8134 8031 8186
rect 8043 8134 8095 8186
rect 14720 8134 14772 8186
rect 14784 8134 14836 8186
rect 14848 8134 14900 8186
rect 14912 8134 14964 8186
rect 4416 7590 4468 7642
rect 4480 7590 4532 7642
rect 4544 7590 4596 7642
rect 4608 7590 4660 7642
rect 11286 7590 11338 7642
rect 11350 7590 11402 7642
rect 11414 7590 11466 7642
rect 11478 7590 11530 7642
rect 18155 7590 18207 7642
rect 18219 7590 18271 7642
rect 18283 7590 18335 7642
rect 18347 7590 18399 7642
rect 7851 7046 7903 7098
rect 7915 7046 7967 7098
rect 7979 7046 8031 7098
rect 8043 7046 8095 7098
rect 14720 7046 14772 7098
rect 14784 7046 14836 7098
rect 14848 7046 14900 7098
rect 14912 7046 14964 7098
rect 4416 6502 4468 6554
rect 4480 6502 4532 6554
rect 4544 6502 4596 6554
rect 4608 6502 4660 6554
rect 11286 6502 11338 6554
rect 11350 6502 11402 6554
rect 11414 6502 11466 6554
rect 11478 6502 11530 6554
rect 18155 6502 18207 6554
rect 18219 6502 18271 6554
rect 18283 6502 18335 6554
rect 18347 6502 18399 6554
rect 7851 5958 7903 6010
rect 7915 5958 7967 6010
rect 7979 5958 8031 6010
rect 8043 5958 8095 6010
rect 14720 5958 14772 6010
rect 14784 5958 14836 6010
rect 14848 5958 14900 6010
rect 14912 5958 14964 6010
rect 4416 5414 4468 5466
rect 4480 5414 4532 5466
rect 4544 5414 4596 5466
rect 4608 5414 4660 5466
rect 11286 5414 11338 5466
rect 11350 5414 11402 5466
rect 11414 5414 11466 5466
rect 11478 5414 11530 5466
rect 18155 5414 18207 5466
rect 18219 5414 18271 5466
rect 18283 5414 18335 5466
rect 18347 5414 18399 5466
rect 7851 4870 7903 4922
rect 7915 4870 7967 4922
rect 7979 4870 8031 4922
rect 8043 4870 8095 4922
rect 14720 4870 14772 4922
rect 14784 4870 14836 4922
rect 14848 4870 14900 4922
rect 14912 4870 14964 4922
rect 4416 4326 4468 4378
rect 4480 4326 4532 4378
rect 4544 4326 4596 4378
rect 4608 4326 4660 4378
rect 11286 4326 11338 4378
rect 11350 4326 11402 4378
rect 11414 4326 11466 4378
rect 11478 4326 11530 4378
rect 18155 4326 18207 4378
rect 18219 4326 18271 4378
rect 18283 4326 18335 4378
rect 18347 4326 18399 4378
rect 9220 4088 9272 4140
rect 11612 4088 11664 4140
rect 6276 4020 6328 4072
rect 11704 4020 11756 4072
rect 7851 3782 7903 3834
rect 7915 3782 7967 3834
rect 7979 3782 8031 3834
rect 8043 3782 8095 3834
rect 14720 3782 14772 3834
rect 14784 3782 14836 3834
rect 14848 3782 14900 3834
rect 14912 3782 14964 3834
rect 572 3476 624 3528
rect 1492 3476 1544 3528
rect 16580 3476 16632 3528
rect 17868 3476 17920 3528
rect 4416 3238 4468 3290
rect 4480 3238 4532 3290
rect 4544 3238 4596 3290
rect 4608 3238 4660 3290
rect 11286 3238 11338 3290
rect 11350 3238 11402 3290
rect 11414 3238 11466 3290
rect 11478 3238 11530 3290
rect 18155 3238 18207 3290
rect 18219 3238 18271 3290
rect 18283 3238 18335 3290
rect 18347 3238 18399 3290
rect 7851 2694 7903 2746
rect 7915 2694 7967 2746
rect 7979 2694 8031 2746
rect 8043 2694 8095 2746
rect 14720 2694 14772 2746
rect 14784 2694 14836 2746
rect 14848 2694 14900 2746
rect 14912 2694 14964 2746
rect 4416 2150 4468 2202
rect 4480 2150 4532 2202
rect 4544 2150 4596 2202
rect 4608 2150 4660 2202
rect 11286 2150 11338 2202
rect 11350 2150 11402 2202
rect 11414 2150 11466 2202
rect 11478 2150 11530 2202
rect 18155 2150 18207 2202
rect 18219 2150 18271 2202
rect 18283 2150 18335 2202
rect 18347 2150 18399 2202
<< metal2 >>
rect 2042 24202 2098 25002
rect 4802 24202 4858 25002
rect 7746 24202 7802 25002
rect 10690 24202 10746 25002
rect 13450 24202 13506 25002
rect 16394 24202 16450 25002
rect 19338 24202 19394 25002
rect 22098 24202 22154 25002
rect 1582 22128 1638 22137
rect 1582 22063 1638 22072
rect 1596 21078 1624 22063
rect 2056 21434 2084 24202
rect 4252 22092 4304 22098
rect 4252 22034 4304 22040
rect 3148 21480 3200 21486
rect 2056 21406 2268 21434
rect 3148 21422 3200 21428
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 2044 21344 2096 21350
rect 2044 21286 2096 21292
rect 1584 21072 1636 21078
rect 1584 21014 1636 21020
rect 1492 20460 1544 20466
rect 1492 20402 1544 20408
rect 1504 19854 1532 20402
rect 1596 20398 1624 21014
rect 2056 21010 2084 21286
rect 2240 21146 2268 21406
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 2044 21004 2096 21010
rect 2044 20946 2096 20952
rect 1584 20392 1636 20398
rect 1584 20334 1636 20340
rect 1596 19922 1624 20334
rect 1584 19916 1636 19922
rect 1584 19858 1636 19864
rect 1492 19848 1544 19854
rect 1492 19790 1544 19796
rect 1504 3534 1532 19790
rect 1768 19168 1820 19174
rect 1768 19110 1820 19116
rect 1780 18834 1808 19110
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 2056 18426 2084 20946
rect 2136 20936 2188 20942
rect 2136 20878 2188 20884
rect 2148 19990 2176 20878
rect 2136 19984 2188 19990
rect 2136 19926 2188 19932
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 2240 18290 2268 21082
rect 2320 20936 2372 20942
rect 2320 20878 2372 20884
rect 2332 20534 2360 20878
rect 2320 20528 2372 20534
rect 2320 20470 2372 20476
rect 2596 20256 2648 20262
rect 2596 20198 2648 20204
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2332 18834 2360 19110
rect 2608 18834 2636 20198
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2596 18828 2648 18834
rect 2596 18770 2648 18776
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2516 17814 2544 18158
rect 2504 17808 2556 17814
rect 2504 17750 2556 17756
rect 2516 17542 2544 17750
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 1596 17202 1624 17478
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 2700 5001 2728 18566
rect 3160 18222 3188 21422
rect 3344 21146 3372 21422
rect 4068 21344 4120 21350
rect 4068 21286 4120 21292
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 4080 21010 4108 21286
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 4264 20806 4292 22034
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4390 21788 4686 21808
rect 4446 21786 4470 21788
rect 4526 21786 4550 21788
rect 4606 21786 4630 21788
rect 4468 21734 4470 21786
rect 4532 21734 4544 21786
rect 4606 21734 4608 21786
rect 4446 21732 4470 21734
rect 4526 21732 4550 21734
rect 4606 21732 4630 21734
rect 4390 21712 4686 21732
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 4390 20700 4686 20720
rect 4446 20698 4470 20700
rect 4526 20698 4550 20700
rect 4606 20698 4630 20700
rect 4468 20646 4470 20698
rect 4532 20646 4544 20698
rect 4606 20646 4608 20698
rect 4446 20644 4470 20646
rect 4526 20644 4550 20646
rect 4606 20644 4630 20646
rect 4390 20624 4686 20644
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 3608 20392 3660 20398
rect 3608 20334 3660 20340
rect 3620 20058 3648 20334
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 4080 19922 4108 20198
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 4264 19310 4292 20470
rect 4724 20398 4752 21830
rect 4816 21690 4844 24202
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 7760 20942 7788 24202
rect 10704 24154 10732 24202
rect 10704 24126 10916 24154
rect 7825 22332 8121 22352
rect 7881 22330 7905 22332
rect 7961 22330 7985 22332
rect 8041 22330 8065 22332
rect 7903 22278 7905 22330
rect 7967 22278 7979 22330
rect 8041 22278 8043 22330
rect 7881 22276 7905 22278
rect 7961 22276 7985 22278
rect 8041 22276 8065 22278
rect 7825 22256 8121 22276
rect 7825 21244 8121 21264
rect 7881 21242 7905 21244
rect 7961 21242 7985 21244
rect 8041 21242 8065 21244
rect 7903 21190 7905 21242
rect 7967 21190 7979 21242
rect 8041 21190 8043 21242
rect 7881 21188 7905 21190
rect 7961 21188 7985 21190
rect 8041 21188 8065 21190
rect 7825 21168 8121 21188
rect 7748 20936 7800 20942
rect 7748 20878 7800 20884
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 7825 20156 8121 20176
rect 7881 20154 7905 20156
rect 7961 20154 7985 20156
rect 8041 20154 8065 20156
rect 7903 20102 7905 20154
rect 7967 20102 7979 20154
rect 8041 20102 8043 20154
rect 7881 20100 7905 20102
rect 7961 20100 7985 20102
rect 8041 20100 8065 20102
rect 7825 20080 8121 20100
rect 4390 19612 4686 19632
rect 4446 19610 4470 19612
rect 4526 19610 4550 19612
rect 4606 19610 4630 19612
rect 4468 19558 4470 19610
rect 4532 19558 4544 19610
rect 4606 19558 4608 19610
rect 4446 19556 4470 19558
rect 4526 19556 4550 19558
rect 4606 19556 4630 19558
rect 4390 19536 4686 19556
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 2792 17785 2820 18158
rect 2778 17776 2834 17785
rect 2778 17711 2780 17720
rect 2832 17711 2834 17720
rect 2780 17682 2832 17688
rect 3068 17678 3096 18158
rect 2872 17672 2924 17678
rect 2792 17620 2872 17626
rect 2792 17614 2924 17620
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 2792 17598 2912 17614
rect 2686 4992 2742 5001
rect 2686 4927 2742 4936
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 584 800 612 3470
rect 2792 898 2820 17598
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2884 17134 2912 17478
rect 4172 17270 4200 18158
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 4264 17066 4292 18566
rect 4390 18524 4686 18544
rect 4446 18522 4470 18524
rect 4526 18522 4550 18524
rect 4606 18522 4630 18524
rect 4468 18470 4470 18522
rect 4532 18470 4544 18522
rect 4606 18470 4608 18522
rect 4446 18468 4470 18470
rect 4526 18468 4550 18470
rect 4606 18468 4630 18470
rect 4390 18448 4686 18468
rect 4724 17746 4752 19110
rect 6472 18970 6500 19246
rect 7825 19068 8121 19088
rect 7881 19066 7905 19068
rect 7961 19066 7985 19068
rect 8041 19066 8065 19068
rect 7903 19014 7905 19066
rect 7967 19014 7979 19066
rect 8041 19014 8043 19066
rect 7881 19012 7905 19014
rect 7961 19012 7985 19014
rect 8041 19012 8065 19014
rect 7825 18992 8121 19012
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4390 17436 4686 17456
rect 4446 17434 4470 17436
rect 4526 17434 4550 17436
rect 4606 17434 4630 17436
rect 4468 17382 4470 17434
rect 4532 17382 4544 17434
rect 4606 17382 4608 17434
rect 4446 17380 4470 17382
rect 4526 17380 4550 17382
rect 4606 17380 4630 17382
rect 4390 17360 4686 17380
rect 5184 17338 5212 18770
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3988 16658 4016 16934
rect 5276 16794 5304 18770
rect 7825 17980 8121 18000
rect 7881 17978 7905 17980
rect 7961 17978 7985 17980
rect 8041 17978 8065 17980
rect 7903 17926 7905 17978
rect 7967 17926 7979 17978
rect 8041 17926 8043 17978
rect 7881 17924 7905 17926
rect 7961 17924 7985 17926
rect 8041 17924 8065 17926
rect 7825 17904 8121 17924
rect 7825 16892 8121 16912
rect 7881 16890 7905 16892
rect 7961 16890 7985 16892
rect 8041 16890 8065 16892
rect 7903 16838 7905 16890
rect 7967 16838 7979 16890
rect 8041 16838 8043 16890
rect 7881 16836 7905 16838
rect 7961 16836 7985 16838
rect 8041 16836 8065 16838
rect 7825 16816 8121 16836
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 4390 16348 4686 16368
rect 4446 16346 4470 16348
rect 4526 16346 4550 16348
rect 4606 16346 4630 16348
rect 4468 16294 4470 16346
rect 4532 16294 4544 16346
rect 4606 16294 4608 16346
rect 4446 16292 4470 16294
rect 4526 16292 4550 16294
rect 4606 16292 4630 16294
rect 4390 16272 4686 16292
rect 7825 15804 8121 15824
rect 7881 15802 7905 15804
rect 7961 15802 7985 15804
rect 8041 15802 8065 15804
rect 7903 15750 7905 15802
rect 7967 15750 7979 15802
rect 8041 15750 8043 15802
rect 7881 15748 7905 15750
rect 7961 15748 7985 15750
rect 8041 15748 8065 15750
rect 7825 15728 8121 15748
rect 4390 15260 4686 15280
rect 4446 15258 4470 15260
rect 4526 15258 4550 15260
rect 4606 15258 4630 15260
rect 4468 15206 4470 15258
rect 4532 15206 4544 15258
rect 4606 15206 4608 15258
rect 4446 15204 4470 15206
rect 4526 15204 4550 15206
rect 4606 15204 4630 15206
rect 4390 15184 4686 15204
rect 7825 14716 8121 14736
rect 7881 14714 7905 14716
rect 7961 14714 7985 14716
rect 8041 14714 8065 14716
rect 7903 14662 7905 14714
rect 7967 14662 7979 14714
rect 8041 14662 8043 14714
rect 7881 14660 7905 14662
rect 7961 14660 7985 14662
rect 8041 14660 8065 14662
rect 7825 14640 8121 14660
rect 4390 14172 4686 14192
rect 4446 14170 4470 14172
rect 4526 14170 4550 14172
rect 4606 14170 4630 14172
rect 4468 14118 4470 14170
rect 4532 14118 4544 14170
rect 4606 14118 4608 14170
rect 4446 14116 4470 14118
rect 4526 14116 4550 14118
rect 4606 14116 4630 14118
rect 4390 14096 4686 14116
rect 3422 13696 3478 13705
rect 3422 13631 3478 13640
rect 3436 12646 3464 13631
rect 7825 13628 8121 13648
rect 7881 13626 7905 13628
rect 7961 13626 7985 13628
rect 8041 13626 8065 13628
rect 7903 13574 7905 13626
rect 7967 13574 7979 13626
rect 8041 13574 8043 13626
rect 7881 13572 7905 13574
rect 7961 13572 7985 13574
rect 8041 13572 8065 13574
rect 7825 13552 8121 13572
rect 4390 13084 4686 13104
rect 4446 13082 4470 13084
rect 4526 13082 4550 13084
rect 4606 13082 4630 13084
rect 4468 13030 4470 13082
rect 4532 13030 4544 13082
rect 4606 13030 4608 13082
rect 4446 13028 4470 13030
rect 4526 13028 4550 13030
rect 4606 13028 4630 13030
rect 4390 13008 4686 13028
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 7825 12540 8121 12560
rect 7881 12538 7905 12540
rect 7961 12538 7985 12540
rect 8041 12538 8065 12540
rect 7903 12486 7905 12538
rect 7967 12486 7979 12538
rect 8041 12486 8043 12538
rect 7881 12484 7905 12486
rect 7961 12484 7985 12486
rect 8041 12484 8065 12486
rect 7825 12464 8121 12484
rect 4390 11996 4686 12016
rect 4446 11994 4470 11996
rect 4526 11994 4550 11996
rect 4606 11994 4630 11996
rect 4468 11942 4470 11994
rect 4532 11942 4544 11994
rect 4606 11942 4608 11994
rect 4446 11940 4470 11942
rect 4526 11940 4550 11942
rect 4606 11940 4630 11942
rect 4390 11920 4686 11940
rect 7825 11452 8121 11472
rect 7881 11450 7905 11452
rect 7961 11450 7985 11452
rect 8041 11450 8065 11452
rect 7903 11398 7905 11450
rect 7967 11398 7979 11450
rect 8041 11398 8043 11450
rect 7881 11396 7905 11398
rect 7961 11396 7985 11398
rect 8041 11396 8065 11398
rect 7825 11376 8121 11396
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 4390 10908 4686 10928
rect 4446 10906 4470 10908
rect 4526 10906 4550 10908
rect 4606 10906 4630 10908
rect 4468 10854 4470 10906
rect 4532 10854 4544 10906
rect 4606 10854 4608 10906
rect 4446 10852 4470 10854
rect 4526 10852 4550 10854
rect 4606 10852 4630 10854
rect 4390 10832 4686 10852
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 7825 10364 8121 10384
rect 7881 10362 7905 10364
rect 7961 10362 7985 10364
rect 8041 10362 8065 10364
rect 7903 10310 7905 10362
rect 7967 10310 7979 10362
rect 8041 10310 8043 10362
rect 7881 10308 7905 10310
rect 7961 10308 7985 10310
rect 8041 10308 8065 10310
rect 7825 10288 8121 10308
rect 10244 10130 10272 10474
rect 10612 10198 10640 10610
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 4390 9820 4686 9840
rect 4446 9818 4470 9820
rect 4526 9818 4550 9820
rect 4606 9818 4630 9820
rect 4468 9766 4470 9818
rect 4532 9766 4544 9818
rect 4606 9766 4608 9818
rect 4446 9764 4470 9766
rect 4526 9764 4550 9766
rect 4606 9764 4630 9766
rect 4390 9744 4686 9764
rect 10244 9518 10272 10066
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 4080 9353 4108 9454
rect 4066 9344 4122 9353
rect 4066 9279 4122 9288
rect 7825 9276 8121 9296
rect 7881 9274 7905 9276
rect 7961 9274 7985 9276
rect 8041 9274 8065 9276
rect 7903 9222 7905 9274
rect 7967 9222 7979 9274
rect 8041 9222 8043 9274
rect 7881 9220 7905 9222
rect 7961 9220 7985 9222
rect 8041 9220 8065 9222
rect 7825 9200 8121 9220
rect 10796 9042 10824 11018
rect 10888 10606 10916 24126
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 11260 21788 11556 21808
rect 11316 21786 11340 21788
rect 11396 21786 11420 21788
rect 11476 21786 11500 21788
rect 11338 21734 11340 21786
rect 11402 21734 11414 21786
rect 11476 21734 11478 21786
rect 11316 21732 11340 21734
rect 11396 21732 11420 21734
rect 11476 21732 11500 21734
rect 11260 21712 11556 21732
rect 13004 21418 13032 21830
rect 13084 21480 13136 21486
rect 13084 21422 13136 21428
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 13096 21146 13124 21422
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 12440 21072 12492 21078
rect 13188 21026 13216 22034
rect 13464 21690 13492 24202
rect 14694 22332 14990 22352
rect 14750 22330 14774 22332
rect 14830 22330 14854 22332
rect 14910 22330 14934 22332
rect 14772 22278 14774 22330
rect 14836 22278 14848 22330
rect 14910 22278 14912 22330
rect 14750 22276 14774 22278
rect 14830 22276 14854 22278
rect 14910 22276 14934 22278
rect 14694 22256 14990 22276
rect 14556 22024 14608 22030
rect 14556 21966 14608 21972
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 12440 21014 12492 21020
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 11260 20700 11556 20720
rect 11316 20698 11340 20700
rect 11396 20698 11420 20700
rect 11476 20698 11500 20700
rect 11338 20646 11340 20698
rect 11402 20646 11414 20698
rect 11476 20646 11478 20698
rect 11316 20644 11340 20646
rect 11396 20644 11420 20646
rect 11476 20644 11500 20646
rect 11260 20624 11556 20644
rect 11900 20058 11928 20946
rect 11888 20052 11940 20058
rect 11888 19994 11940 20000
rect 12452 19922 12480 21014
rect 12716 21004 12768 21010
rect 12716 20946 12768 20952
rect 13096 20998 13216 21026
rect 13360 21004 13412 21010
rect 12728 20602 12756 20946
rect 13096 20874 13124 20998
rect 13360 20946 13412 20952
rect 13084 20868 13136 20874
rect 13084 20810 13136 20816
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12728 19922 12756 20538
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 11260 19612 11556 19632
rect 11316 19610 11340 19612
rect 11396 19610 11420 19612
rect 11476 19610 11500 19612
rect 11338 19558 11340 19610
rect 11402 19558 11414 19610
rect 11476 19558 11478 19610
rect 11316 19556 11340 19558
rect 11396 19556 11420 19558
rect 11476 19556 11500 19558
rect 11260 19536 11556 19556
rect 12820 19310 12848 20742
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 13004 19990 13032 20402
rect 13096 20398 13124 20810
rect 13372 20466 13400 20946
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 12992 19984 13044 19990
rect 12992 19926 13044 19932
rect 13832 19922 13860 21830
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 11260 18524 11556 18544
rect 11316 18522 11340 18524
rect 11396 18522 11420 18524
rect 11476 18522 11500 18524
rect 11338 18470 11340 18522
rect 11402 18470 11414 18522
rect 11476 18470 11478 18522
rect 11316 18468 11340 18470
rect 11396 18468 11420 18470
rect 11476 18468 11500 18470
rect 11260 18448 11556 18468
rect 11260 17436 11556 17456
rect 11316 17434 11340 17436
rect 11396 17434 11420 17436
rect 11476 17434 11500 17436
rect 11338 17382 11340 17434
rect 11402 17382 11414 17434
rect 11476 17382 11478 17434
rect 11316 17380 11340 17382
rect 11396 17380 11420 17382
rect 11476 17380 11500 17382
rect 11260 17360 11556 17380
rect 11260 16348 11556 16368
rect 11316 16346 11340 16348
rect 11396 16346 11420 16348
rect 11476 16346 11500 16348
rect 11338 16294 11340 16346
rect 11402 16294 11414 16346
rect 11476 16294 11478 16346
rect 11316 16292 11340 16294
rect 11396 16292 11420 16294
rect 11476 16292 11500 16294
rect 11260 16272 11556 16292
rect 11260 15260 11556 15280
rect 11316 15258 11340 15260
rect 11396 15258 11420 15260
rect 11476 15258 11500 15260
rect 11338 15206 11340 15258
rect 11402 15206 11414 15258
rect 11476 15206 11478 15258
rect 11316 15204 11340 15206
rect 11396 15204 11420 15206
rect 11476 15204 11500 15206
rect 11260 15184 11556 15204
rect 11260 14172 11556 14192
rect 11316 14170 11340 14172
rect 11396 14170 11420 14172
rect 11476 14170 11500 14172
rect 11338 14118 11340 14170
rect 11402 14118 11414 14170
rect 11476 14118 11478 14170
rect 11316 14116 11340 14118
rect 11396 14116 11420 14118
rect 11476 14116 11500 14118
rect 11260 14096 11556 14116
rect 11260 13084 11556 13104
rect 11316 13082 11340 13084
rect 11396 13082 11420 13084
rect 11476 13082 11500 13084
rect 11338 13030 11340 13082
rect 11402 13030 11414 13082
rect 11476 13030 11478 13082
rect 11316 13028 11340 13030
rect 11396 13028 11420 13030
rect 11476 13028 11500 13030
rect 11260 13008 11556 13028
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 11260 11996 11556 12016
rect 11316 11994 11340 11996
rect 11396 11994 11420 11996
rect 11476 11994 11500 11996
rect 11338 11942 11340 11994
rect 11402 11942 11414 11994
rect 11476 11942 11478 11994
rect 11316 11940 11340 11942
rect 11396 11940 11420 11942
rect 11476 11940 11500 11942
rect 11260 11920 11556 11940
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 11072 10674 11100 11154
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 11260 10908 11556 10928
rect 11316 10906 11340 10908
rect 11396 10906 11420 10908
rect 11476 10906 11500 10908
rect 11338 10854 11340 10906
rect 11402 10854 11414 10906
rect 11476 10854 11478 10906
rect 11316 10852 11340 10854
rect 11396 10852 11420 10854
rect 11476 10852 11500 10854
rect 11260 10832 11556 10852
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10888 10062 10916 10542
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10888 9518 10916 9998
rect 11260 9820 11556 9840
rect 11316 9818 11340 9820
rect 11396 9818 11420 9820
rect 11476 9818 11500 9820
rect 11338 9766 11340 9818
rect 11402 9766 11414 9818
rect 11476 9766 11478 9818
rect 11316 9764 11340 9766
rect 11396 9764 11420 9766
rect 11476 9764 11500 9766
rect 11260 9744 11556 9764
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 9042 10916 9318
rect 11624 9110 11652 10066
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 4390 8732 4686 8752
rect 4446 8730 4470 8732
rect 4526 8730 4550 8732
rect 4606 8730 4630 8732
rect 4468 8678 4470 8730
rect 4532 8678 4544 8730
rect 4606 8678 4608 8730
rect 4446 8676 4470 8678
rect 4526 8676 4550 8678
rect 4606 8676 4630 8678
rect 4390 8656 4686 8676
rect 11164 8634 11192 8978
rect 11260 8732 11556 8752
rect 11316 8730 11340 8732
rect 11396 8730 11420 8732
rect 11476 8730 11500 8732
rect 11338 8678 11340 8730
rect 11402 8678 11414 8730
rect 11476 8678 11478 8730
rect 11316 8676 11340 8678
rect 11396 8676 11420 8678
rect 11476 8676 11500 8678
rect 11260 8656 11556 8676
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 7825 8188 8121 8208
rect 7881 8186 7905 8188
rect 7961 8186 7985 8188
rect 8041 8186 8065 8188
rect 7903 8134 7905 8186
rect 7967 8134 7979 8186
rect 8041 8134 8043 8186
rect 7881 8132 7905 8134
rect 7961 8132 7985 8134
rect 8041 8132 8065 8134
rect 7825 8112 8121 8132
rect 4390 7644 4686 7664
rect 4446 7642 4470 7644
rect 4526 7642 4550 7644
rect 4606 7642 4630 7644
rect 4468 7590 4470 7642
rect 4532 7590 4544 7642
rect 4606 7590 4608 7642
rect 4446 7588 4470 7590
rect 4526 7588 4550 7590
rect 4606 7588 4630 7590
rect 4390 7568 4686 7588
rect 11260 7644 11556 7664
rect 11316 7642 11340 7644
rect 11396 7642 11420 7644
rect 11476 7642 11500 7644
rect 11338 7590 11340 7642
rect 11402 7590 11414 7642
rect 11476 7590 11478 7642
rect 11316 7588 11340 7590
rect 11396 7588 11420 7590
rect 11476 7588 11500 7590
rect 11260 7568 11556 7588
rect 7825 7100 8121 7120
rect 7881 7098 7905 7100
rect 7961 7098 7985 7100
rect 8041 7098 8065 7100
rect 7903 7046 7905 7098
rect 7967 7046 7979 7098
rect 8041 7046 8043 7098
rect 7881 7044 7905 7046
rect 7961 7044 7985 7046
rect 8041 7044 8065 7046
rect 7825 7024 8121 7044
rect 4390 6556 4686 6576
rect 4446 6554 4470 6556
rect 4526 6554 4550 6556
rect 4606 6554 4630 6556
rect 4468 6502 4470 6554
rect 4532 6502 4544 6554
rect 4606 6502 4608 6554
rect 4446 6500 4470 6502
rect 4526 6500 4550 6502
rect 4606 6500 4630 6502
rect 4390 6480 4686 6500
rect 11260 6556 11556 6576
rect 11316 6554 11340 6556
rect 11396 6554 11420 6556
rect 11476 6554 11500 6556
rect 11338 6502 11340 6554
rect 11402 6502 11414 6554
rect 11476 6502 11478 6554
rect 11316 6500 11340 6502
rect 11396 6500 11420 6502
rect 11476 6500 11500 6502
rect 11260 6480 11556 6500
rect 7825 6012 8121 6032
rect 7881 6010 7905 6012
rect 7961 6010 7985 6012
rect 8041 6010 8065 6012
rect 7903 5958 7905 6010
rect 7967 5958 7979 6010
rect 8041 5958 8043 6010
rect 7881 5956 7905 5958
rect 7961 5956 7985 5958
rect 8041 5956 8065 5958
rect 7825 5936 8121 5956
rect 4390 5468 4686 5488
rect 4446 5466 4470 5468
rect 4526 5466 4550 5468
rect 4606 5466 4630 5468
rect 4468 5414 4470 5466
rect 4532 5414 4544 5466
rect 4606 5414 4608 5466
rect 4446 5412 4470 5414
rect 4526 5412 4550 5414
rect 4606 5412 4630 5414
rect 4390 5392 4686 5412
rect 11260 5468 11556 5488
rect 11316 5466 11340 5468
rect 11396 5466 11420 5468
rect 11476 5466 11500 5468
rect 11338 5414 11340 5466
rect 11402 5414 11414 5466
rect 11476 5414 11478 5466
rect 11316 5412 11340 5414
rect 11396 5412 11420 5414
rect 11476 5412 11500 5414
rect 11260 5392 11556 5412
rect 7825 4924 8121 4944
rect 7881 4922 7905 4924
rect 7961 4922 7985 4924
rect 8041 4922 8065 4924
rect 7903 4870 7905 4922
rect 7967 4870 7979 4922
rect 8041 4870 8043 4922
rect 7881 4868 7905 4870
rect 7961 4868 7985 4870
rect 8041 4868 8065 4870
rect 7825 4848 8121 4868
rect 4390 4380 4686 4400
rect 4446 4378 4470 4380
rect 4526 4378 4550 4380
rect 4606 4378 4630 4380
rect 4468 4326 4470 4378
rect 4532 4326 4544 4378
rect 4606 4326 4608 4378
rect 4446 4324 4470 4326
rect 4526 4324 4550 4326
rect 4606 4324 4630 4326
rect 4390 4304 4686 4324
rect 11260 4380 11556 4400
rect 11316 4378 11340 4380
rect 11396 4378 11420 4380
rect 11476 4378 11500 4380
rect 11338 4326 11340 4378
rect 11402 4326 11414 4378
rect 11476 4326 11478 4378
rect 11316 4324 11340 4326
rect 11396 4324 11420 4326
rect 11476 4324 11500 4326
rect 11260 4304 11556 4324
rect 11624 4146 11652 9046
rect 11808 8974 11836 10610
rect 12820 10606 12848 10950
rect 13372 10606 13400 10950
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 12912 10198 12940 10542
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12360 10010 12388 10066
rect 12268 9982 12388 10010
rect 12268 9518 12296 9982
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 4390 3292 4686 3312
rect 4446 3290 4470 3292
rect 4526 3290 4550 3292
rect 4606 3290 4630 3292
rect 4468 3238 4470 3290
rect 4532 3238 4544 3290
rect 4606 3238 4608 3290
rect 4446 3236 4470 3238
rect 4526 3236 4550 3238
rect 4606 3236 4630 3238
rect 4390 3216 4686 3236
rect 4390 2204 4686 2224
rect 4446 2202 4470 2204
rect 4526 2202 4550 2204
rect 4606 2202 4630 2204
rect 4468 2150 4470 2202
rect 4532 2150 4544 2202
rect 4606 2150 4608 2202
rect 4446 2148 4470 2150
rect 4526 2148 4550 2150
rect 4606 2148 4630 2150
rect 4390 2128 4686 2148
rect 2792 870 3372 898
rect 3344 800 3372 870
rect 6288 800 6316 4014
rect 7825 3836 8121 3856
rect 7881 3834 7905 3836
rect 7961 3834 7985 3836
rect 8041 3834 8065 3836
rect 7903 3782 7905 3834
rect 7967 3782 7979 3834
rect 8041 3782 8043 3834
rect 7881 3780 7905 3782
rect 7961 3780 7985 3782
rect 8041 3780 8065 3782
rect 7825 3760 8121 3780
rect 7825 2748 8121 2768
rect 7881 2746 7905 2748
rect 7961 2746 7985 2748
rect 8041 2746 8065 2748
rect 7903 2694 7905 2746
rect 7967 2694 7979 2746
rect 8041 2694 8043 2746
rect 7881 2692 7905 2694
rect 7961 2692 7985 2694
rect 8041 2692 8065 2694
rect 7825 2672 8121 2692
rect 9232 800 9260 4082
rect 11716 4078 11744 8842
rect 11808 8430 11836 8910
rect 12268 8906 12296 9454
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 12360 9110 12388 9386
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 13280 9042 13308 9386
rect 13464 9042 13492 11154
rect 13924 10742 13952 12582
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13924 10130 13952 10678
rect 14108 10674 14136 21354
rect 14568 20602 14596 21966
rect 14694 21244 14990 21264
rect 14750 21242 14774 21244
rect 14830 21242 14854 21244
rect 14910 21242 14934 21244
rect 14772 21190 14774 21242
rect 14836 21190 14848 21242
rect 14910 21190 14912 21242
rect 14750 21188 14774 21190
rect 14830 21188 14854 21190
rect 14910 21188 14934 21190
rect 14694 21168 14990 21188
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 14694 20156 14990 20176
rect 14750 20154 14774 20156
rect 14830 20154 14854 20156
rect 14910 20154 14934 20156
rect 14772 20102 14774 20154
rect 14836 20102 14848 20154
rect 14910 20102 14912 20154
rect 14750 20100 14774 20102
rect 14830 20100 14854 20102
rect 14910 20100 14934 20102
rect 14694 20080 14990 20100
rect 14694 19068 14990 19088
rect 14750 19066 14774 19068
rect 14830 19066 14854 19068
rect 14910 19066 14934 19068
rect 14772 19014 14774 19066
rect 14836 19014 14848 19066
rect 14910 19014 14912 19066
rect 14750 19012 14774 19014
rect 14830 19012 14854 19014
rect 14910 19012 14934 19014
rect 14694 18992 14990 19012
rect 14694 17980 14990 18000
rect 14750 17978 14774 17980
rect 14830 17978 14854 17980
rect 14910 17978 14934 17980
rect 14772 17926 14774 17978
rect 14836 17926 14848 17978
rect 14910 17926 14912 17978
rect 14750 17924 14774 17926
rect 14830 17924 14854 17926
rect 14910 17924 14934 17926
rect 14694 17904 14990 17924
rect 14694 16892 14990 16912
rect 14750 16890 14774 16892
rect 14830 16890 14854 16892
rect 14910 16890 14934 16892
rect 14772 16838 14774 16890
rect 14836 16838 14848 16890
rect 14910 16838 14912 16890
rect 14750 16836 14774 16838
rect 14830 16836 14854 16838
rect 14910 16836 14934 16838
rect 14694 16816 14990 16836
rect 14694 15804 14990 15824
rect 14750 15802 14774 15804
rect 14830 15802 14854 15804
rect 14910 15802 14934 15804
rect 14772 15750 14774 15802
rect 14836 15750 14848 15802
rect 14910 15750 14912 15802
rect 14750 15748 14774 15750
rect 14830 15748 14854 15750
rect 14910 15748 14934 15750
rect 14694 15728 14990 15748
rect 14694 14716 14990 14736
rect 14750 14714 14774 14716
rect 14830 14714 14854 14716
rect 14910 14714 14934 14716
rect 14772 14662 14774 14714
rect 14836 14662 14848 14714
rect 14910 14662 14912 14714
rect 14750 14660 14774 14662
rect 14830 14660 14854 14662
rect 14910 14660 14934 14662
rect 14694 14640 14990 14660
rect 14694 13628 14990 13648
rect 14750 13626 14774 13628
rect 14830 13626 14854 13628
rect 14910 13626 14934 13628
rect 14772 13574 14774 13626
rect 14836 13574 14848 13626
rect 14910 13574 14912 13626
rect 14750 13572 14774 13574
rect 14830 13572 14854 13574
rect 14910 13572 14934 13574
rect 14694 13552 14990 13572
rect 14694 12540 14990 12560
rect 14750 12538 14774 12540
rect 14830 12538 14854 12540
rect 14910 12538 14934 12540
rect 14772 12486 14774 12538
rect 14836 12486 14848 12538
rect 14910 12486 14912 12538
rect 14750 12484 14774 12486
rect 14830 12484 14854 12486
rect 14910 12484 14934 12486
rect 14694 12464 14990 12484
rect 14694 11452 14990 11472
rect 14750 11450 14774 11452
rect 14830 11450 14854 11452
rect 14910 11450 14934 11452
rect 14772 11398 14774 11450
rect 14836 11398 14848 11450
rect 14910 11398 14912 11450
rect 14750 11396 14774 11398
rect 14830 11396 14854 11398
rect 14910 11396 14934 11398
rect 14694 11376 14990 11396
rect 15212 10810 15240 20402
rect 15304 19174 15332 20946
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15488 20398 15516 20742
rect 16408 20466 16436 24202
rect 18129 21788 18425 21808
rect 18185 21786 18209 21788
rect 18265 21786 18289 21788
rect 18345 21786 18369 21788
rect 18207 21734 18209 21786
rect 18271 21734 18283 21786
rect 18345 21734 18347 21786
rect 18185 21732 18209 21734
rect 18265 21732 18289 21734
rect 18345 21732 18369 21734
rect 18129 21712 18425 21732
rect 19352 21418 19380 24202
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 18129 20700 18425 20720
rect 18185 20698 18209 20700
rect 18265 20698 18289 20700
rect 18345 20698 18369 20700
rect 18207 20646 18209 20698
rect 18271 20646 18283 20698
rect 18345 20646 18347 20698
rect 18185 20644 18209 20646
rect 18265 20644 18289 20646
rect 18345 20644 18369 20646
rect 18129 20624 18425 20644
rect 22112 20466 22140 24202
rect 16396 20460 16448 20466
rect 16396 20402 16448 20408
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 17684 20256 17736 20262
rect 17684 20198 17736 20204
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16776 11354 16804 12242
rect 17696 12186 17724 20198
rect 18432 19961 18460 20402
rect 18418 19952 18474 19961
rect 18418 19887 18474 19896
rect 18129 19612 18425 19632
rect 18185 19610 18209 19612
rect 18265 19610 18289 19612
rect 18345 19610 18369 19612
rect 18207 19558 18209 19610
rect 18271 19558 18283 19610
rect 18345 19558 18347 19610
rect 18185 19556 18209 19558
rect 18265 19556 18289 19558
rect 18345 19556 18369 19558
rect 18129 19536 18425 19556
rect 18129 18524 18425 18544
rect 18185 18522 18209 18524
rect 18265 18522 18289 18524
rect 18345 18522 18369 18524
rect 18207 18470 18209 18522
rect 18271 18470 18283 18522
rect 18345 18470 18347 18522
rect 18185 18468 18209 18470
rect 18265 18468 18289 18470
rect 18345 18468 18369 18470
rect 18129 18448 18425 18468
rect 18129 17436 18425 17456
rect 18185 17434 18209 17436
rect 18265 17434 18289 17436
rect 18345 17434 18369 17436
rect 18207 17382 18209 17434
rect 18271 17382 18283 17434
rect 18345 17382 18347 17434
rect 18185 17380 18209 17382
rect 18265 17380 18289 17382
rect 18345 17380 18369 17382
rect 18129 17360 18425 17380
rect 18129 16348 18425 16368
rect 18185 16346 18209 16348
rect 18265 16346 18289 16348
rect 18345 16346 18369 16348
rect 18207 16294 18209 16346
rect 18271 16294 18283 16346
rect 18345 16294 18347 16346
rect 18185 16292 18209 16294
rect 18265 16292 18289 16294
rect 18345 16292 18369 16294
rect 18129 16272 18425 16292
rect 19522 15600 19578 15609
rect 19522 15535 19578 15544
rect 18129 15260 18425 15280
rect 18185 15258 18209 15260
rect 18265 15258 18289 15260
rect 18345 15258 18369 15260
rect 18207 15206 18209 15258
rect 18271 15206 18283 15258
rect 18345 15206 18347 15258
rect 18185 15204 18209 15206
rect 18265 15204 18289 15206
rect 18345 15204 18369 15206
rect 18129 15184 18425 15204
rect 18129 14172 18425 14192
rect 18185 14170 18209 14172
rect 18265 14170 18289 14172
rect 18345 14170 18369 14172
rect 18207 14118 18209 14170
rect 18271 14118 18283 14170
rect 18345 14118 18347 14170
rect 18185 14116 18209 14118
rect 18265 14116 18289 14118
rect 18345 14116 18369 14118
rect 18129 14096 18425 14116
rect 18129 13084 18425 13104
rect 18185 13082 18209 13084
rect 18265 13082 18289 13084
rect 18345 13082 18369 13084
rect 18207 13030 18209 13082
rect 18271 13030 18283 13082
rect 18345 13030 18347 13082
rect 18185 13028 18209 13030
rect 18265 13028 18289 13030
rect 18345 13028 18369 13030
rect 18129 13008 18425 13028
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 17604 12158 17724 12186
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13924 9518 13952 10066
rect 14108 10062 14136 10610
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14384 10198 14412 10542
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 14694 10364 14990 10384
rect 14750 10362 14774 10364
rect 14830 10362 14854 10364
rect 14910 10362 14934 10364
rect 14772 10310 14774 10362
rect 14836 10310 14848 10362
rect 14910 10310 14912 10362
rect 14750 10308 14774 10310
rect 14830 10308 14854 10310
rect 14910 10308 14934 10310
rect 14694 10288 14990 10308
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 15212 10130 15240 10474
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14108 9518 14136 9998
rect 15108 9988 15160 9994
rect 15108 9930 15160 9936
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14694 9276 14990 9296
rect 14750 9274 14774 9276
rect 14830 9274 14854 9276
rect 14910 9274 14934 9276
rect 14772 9222 14774 9274
rect 14836 9222 14848 9274
rect 14910 9222 14912 9274
rect 14750 9220 14774 9222
rect 14830 9220 14854 9222
rect 14910 9220 14934 9222
rect 14694 9200 14990 9220
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11260 3292 11556 3312
rect 11316 3290 11340 3292
rect 11396 3290 11420 3292
rect 11476 3290 11500 3292
rect 11338 3238 11340 3290
rect 11402 3238 11414 3290
rect 11476 3238 11478 3290
rect 11316 3236 11340 3238
rect 11396 3236 11420 3238
rect 11476 3236 11500 3238
rect 11260 3216 11556 3236
rect 11260 2204 11556 2224
rect 11316 2202 11340 2204
rect 11396 2202 11420 2204
rect 11476 2202 11500 2204
rect 11338 2150 11340 2202
rect 11402 2150 11414 2202
rect 11476 2150 11478 2202
rect 11316 2148 11340 2150
rect 11396 2148 11420 2150
rect 11476 2148 11500 2150
rect 11260 2128 11556 2148
rect 11992 800 12020 8774
rect 14694 8188 14990 8208
rect 14750 8186 14774 8188
rect 14830 8186 14854 8188
rect 14910 8186 14934 8188
rect 14772 8134 14774 8186
rect 14836 8134 14848 8186
rect 14910 8134 14912 8186
rect 14750 8132 14774 8134
rect 14830 8132 14854 8134
rect 14910 8132 14934 8134
rect 14694 8112 14990 8132
rect 14694 7100 14990 7120
rect 14750 7098 14774 7100
rect 14830 7098 14854 7100
rect 14910 7098 14934 7100
rect 14772 7046 14774 7098
rect 14836 7046 14848 7098
rect 14910 7046 14912 7098
rect 14750 7044 14774 7046
rect 14830 7044 14854 7046
rect 14910 7044 14934 7046
rect 14694 7024 14990 7044
rect 14694 6012 14990 6032
rect 14750 6010 14774 6012
rect 14830 6010 14854 6012
rect 14910 6010 14934 6012
rect 14772 5958 14774 6010
rect 14836 5958 14848 6010
rect 14910 5958 14912 6010
rect 14750 5956 14774 5958
rect 14830 5956 14854 5958
rect 14910 5956 14934 5958
rect 14694 5936 14990 5956
rect 14694 4924 14990 4944
rect 14750 4922 14774 4924
rect 14830 4922 14854 4924
rect 14910 4922 14934 4924
rect 14772 4870 14774 4922
rect 14836 4870 14848 4922
rect 14910 4870 14912 4922
rect 14750 4868 14774 4870
rect 14830 4868 14854 4870
rect 14910 4868 14934 4870
rect 14694 4848 14990 4868
rect 14694 3836 14990 3856
rect 14750 3834 14774 3836
rect 14830 3834 14854 3836
rect 14910 3834 14934 3836
rect 14772 3782 14774 3834
rect 14836 3782 14848 3834
rect 14910 3782 14912 3834
rect 14750 3780 14774 3782
rect 14830 3780 14854 3782
rect 14910 3780 14934 3782
rect 14694 3760 14990 3780
rect 14694 2748 14990 2768
rect 14750 2746 14774 2748
rect 14830 2746 14854 2748
rect 14910 2746 14934 2748
rect 14772 2694 14774 2746
rect 14836 2694 14848 2746
rect 14910 2694 14912 2746
rect 14750 2692 14774 2694
rect 14830 2692 14854 2694
rect 14910 2692 14934 2694
rect 14694 2672 14990 2692
rect 15120 2394 15148 9930
rect 15488 9586 15516 10066
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 16592 3534 16620 10406
rect 17604 10130 17632 12158
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17696 11218 17724 12038
rect 18129 11996 18425 12016
rect 18185 11994 18209 11996
rect 18265 11994 18289 11996
rect 18345 11994 18369 11996
rect 18207 11942 18209 11994
rect 18271 11942 18283 11994
rect 18345 11942 18347 11994
rect 18185 11940 18209 11942
rect 18265 11940 18289 11942
rect 18345 11940 18369 11942
rect 18129 11920 18425 11940
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17880 11354 17908 11630
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 18064 10606 18092 11494
rect 19352 11218 19380 12718
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19352 11098 19380 11154
rect 19260 11070 19380 11098
rect 18129 10908 18425 10928
rect 18185 10906 18209 10908
rect 18265 10906 18289 10908
rect 18345 10906 18369 10908
rect 18207 10854 18209 10906
rect 18271 10854 18283 10906
rect 18345 10854 18347 10906
rect 18185 10852 18209 10854
rect 18265 10852 18289 10854
rect 18345 10852 18369 10854
rect 18129 10832 18425 10852
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 19260 10266 19288 11070
rect 19444 10606 19472 12582
rect 19536 12306 19564 15535
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19536 12186 19564 12242
rect 20732 12238 20760 20402
rect 20720 12232 20772 12238
rect 19536 12158 19656 12186
rect 20720 12174 20772 12180
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19536 11150 19564 12038
rect 19628 11694 19656 12158
rect 20732 11694 20760 12174
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 19628 11218 19656 11630
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 19706 11248 19762 11257
rect 19616 11212 19668 11218
rect 19706 11183 19762 11192
rect 19616 11154 19668 11160
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 19720 10062 19748 11183
rect 20456 10606 20484 11494
rect 20732 11218 20760 11630
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 18129 9820 18425 9840
rect 18185 9818 18209 9820
rect 18265 9818 18289 9820
rect 18345 9818 18369 9820
rect 18207 9766 18209 9818
rect 18271 9766 18283 9818
rect 18345 9766 18347 9818
rect 18185 9764 18209 9766
rect 18265 9764 18289 9766
rect 18345 9764 18369 9766
rect 18129 9744 18425 9764
rect 19076 9518 19104 9862
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 19536 8838 19564 9998
rect 19720 8974 19748 9998
rect 19996 9042 20024 10066
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20180 9518 20208 9590
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 18129 8732 18425 8752
rect 18185 8730 18209 8732
rect 18265 8730 18289 8732
rect 18345 8730 18369 8732
rect 18207 8678 18209 8730
rect 18271 8678 18283 8730
rect 18345 8678 18347 8730
rect 18185 8676 18209 8678
rect 18265 8676 18289 8678
rect 18345 8676 18369 8678
rect 18129 8656 18425 8676
rect 19720 8514 19748 8910
rect 19628 8486 19748 8514
rect 19628 8430 19656 8486
rect 19996 8430 20024 8978
rect 20180 8566 20208 9454
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20168 8560 20220 8566
rect 20168 8502 20220 8508
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 18129 7644 18425 7664
rect 18185 7642 18209 7644
rect 18265 7642 18289 7644
rect 18345 7642 18369 7644
rect 18207 7590 18209 7642
rect 18271 7590 18283 7642
rect 18345 7590 18347 7642
rect 18185 7588 18209 7590
rect 18265 7588 18289 7590
rect 18345 7588 18369 7590
rect 18129 7568 18425 7588
rect 19996 7177 20024 8366
rect 19982 7168 20038 7177
rect 19982 7103 20038 7112
rect 18129 6556 18425 6576
rect 18185 6554 18209 6556
rect 18265 6554 18289 6556
rect 18345 6554 18369 6556
rect 18207 6502 18209 6554
rect 18271 6502 18283 6554
rect 18345 6502 18347 6554
rect 18185 6500 18209 6502
rect 18265 6500 18289 6502
rect 18345 6500 18369 6502
rect 18129 6480 18425 6500
rect 18129 5468 18425 5488
rect 18185 5466 18209 5468
rect 18265 5466 18289 5468
rect 18345 5466 18369 5468
rect 18207 5414 18209 5466
rect 18271 5414 18283 5466
rect 18345 5414 18347 5466
rect 18185 5412 18209 5414
rect 18265 5412 18289 5414
rect 18345 5412 18369 5414
rect 18129 5392 18425 5412
rect 18129 4380 18425 4400
rect 18185 4378 18209 4380
rect 18265 4378 18289 4380
rect 18345 4378 18369 4380
rect 18207 4326 18209 4378
rect 18271 4326 18283 4378
rect 18345 4326 18347 4378
rect 18185 4324 18209 4326
rect 18265 4324 18289 4326
rect 18345 4324 18369 4326
rect 18129 4304 18425 4324
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 14936 2366 15148 2394
rect 14936 800 14964 2366
rect 17880 800 17908 3470
rect 18129 3292 18425 3312
rect 18185 3290 18209 3292
rect 18265 3290 18289 3292
rect 18345 3290 18369 3292
rect 18207 3238 18209 3290
rect 18271 3238 18283 3290
rect 18345 3238 18347 3290
rect 18185 3236 18209 3238
rect 18265 3236 18289 3238
rect 18345 3236 18369 3238
rect 18129 3216 18425 3236
rect 20364 2825 20392 9318
rect 20350 2816 20406 2825
rect 20350 2751 20406 2760
rect 18129 2204 18425 2224
rect 18185 2202 18209 2204
rect 18265 2202 18289 2204
rect 18345 2202 18369 2204
rect 18207 2150 18209 2202
rect 18271 2150 18283 2202
rect 18345 2150 18347 2202
rect 18185 2148 18209 2150
rect 18265 2148 18289 2150
rect 18345 2148 18369 2150
rect 18129 2128 18425 2148
rect 20456 898 20484 10406
rect 20456 870 20668 898
rect 20640 800 20668 870
rect 570 0 626 800
rect 3330 0 3386 800
rect 6274 0 6330 800
rect 9218 0 9274 800
rect 11978 0 12034 800
rect 14922 0 14978 800
rect 17866 0 17922 800
rect 20626 0 20682 800
<< via2 >>
rect 1582 22072 1638 22128
rect 4390 21786 4446 21788
rect 4470 21786 4526 21788
rect 4550 21786 4606 21788
rect 4630 21786 4686 21788
rect 4390 21734 4416 21786
rect 4416 21734 4446 21786
rect 4470 21734 4480 21786
rect 4480 21734 4526 21786
rect 4550 21734 4596 21786
rect 4596 21734 4606 21786
rect 4630 21734 4660 21786
rect 4660 21734 4686 21786
rect 4390 21732 4446 21734
rect 4470 21732 4526 21734
rect 4550 21732 4606 21734
rect 4630 21732 4686 21734
rect 4390 20698 4446 20700
rect 4470 20698 4526 20700
rect 4550 20698 4606 20700
rect 4630 20698 4686 20700
rect 4390 20646 4416 20698
rect 4416 20646 4446 20698
rect 4470 20646 4480 20698
rect 4480 20646 4526 20698
rect 4550 20646 4596 20698
rect 4596 20646 4606 20698
rect 4630 20646 4660 20698
rect 4660 20646 4686 20698
rect 4390 20644 4446 20646
rect 4470 20644 4526 20646
rect 4550 20644 4606 20646
rect 4630 20644 4686 20646
rect 7825 22330 7881 22332
rect 7905 22330 7961 22332
rect 7985 22330 8041 22332
rect 8065 22330 8121 22332
rect 7825 22278 7851 22330
rect 7851 22278 7881 22330
rect 7905 22278 7915 22330
rect 7915 22278 7961 22330
rect 7985 22278 8031 22330
rect 8031 22278 8041 22330
rect 8065 22278 8095 22330
rect 8095 22278 8121 22330
rect 7825 22276 7881 22278
rect 7905 22276 7961 22278
rect 7985 22276 8041 22278
rect 8065 22276 8121 22278
rect 7825 21242 7881 21244
rect 7905 21242 7961 21244
rect 7985 21242 8041 21244
rect 8065 21242 8121 21244
rect 7825 21190 7851 21242
rect 7851 21190 7881 21242
rect 7905 21190 7915 21242
rect 7915 21190 7961 21242
rect 7985 21190 8031 21242
rect 8031 21190 8041 21242
rect 8065 21190 8095 21242
rect 8095 21190 8121 21242
rect 7825 21188 7881 21190
rect 7905 21188 7961 21190
rect 7985 21188 8041 21190
rect 8065 21188 8121 21190
rect 7825 20154 7881 20156
rect 7905 20154 7961 20156
rect 7985 20154 8041 20156
rect 8065 20154 8121 20156
rect 7825 20102 7851 20154
rect 7851 20102 7881 20154
rect 7905 20102 7915 20154
rect 7915 20102 7961 20154
rect 7985 20102 8031 20154
rect 8031 20102 8041 20154
rect 8065 20102 8095 20154
rect 8095 20102 8121 20154
rect 7825 20100 7881 20102
rect 7905 20100 7961 20102
rect 7985 20100 8041 20102
rect 8065 20100 8121 20102
rect 4390 19610 4446 19612
rect 4470 19610 4526 19612
rect 4550 19610 4606 19612
rect 4630 19610 4686 19612
rect 4390 19558 4416 19610
rect 4416 19558 4446 19610
rect 4470 19558 4480 19610
rect 4480 19558 4526 19610
rect 4550 19558 4596 19610
rect 4596 19558 4606 19610
rect 4630 19558 4660 19610
rect 4660 19558 4686 19610
rect 4390 19556 4446 19558
rect 4470 19556 4526 19558
rect 4550 19556 4606 19558
rect 4630 19556 4686 19558
rect 2778 17740 2834 17776
rect 2778 17720 2780 17740
rect 2780 17720 2832 17740
rect 2832 17720 2834 17740
rect 2686 4936 2742 4992
rect 4390 18522 4446 18524
rect 4470 18522 4526 18524
rect 4550 18522 4606 18524
rect 4630 18522 4686 18524
rect 4390 18470 4416 18522
rect 4416 18470 4446 18522
rect 4470 18470 4480 18522
rect 4480 18470 4526 18522
rect 4550 18470 4596 18522
rect 4596 18470 4606 18522
rect 4630 18470 4660 18522
rect 4660 18470 4686 18522
rect 4390 18468 4446 18470
rect 4470 18468 4526 18470
rect 4550 18468 4606 18470
rect 4630 18468 4686 18470
rect 7825 19066 7881 19068
rect 7905 19066 7961 19068
rect 7985 19066 8041 19068
rect 8065 19066 8121 19068
rect 7825 19014 7851 19066
rect 7851 19014 7881 19066
rect 7905 19014 7915 19066
rect 7915 19014 7961 19066
rect 7985 19014 8031 19066
rect 8031 19014 8041 19066
rect 8065 19014 8095 19066
rect 8095 19014 8121 19066
rect 7825 19012 7881 19014
rect 7905 19012 7961 19014
rect 7985 19012 8041 19014
rect 8065 19012 8121 19014
rect 4390 17434 4446 17436
rect 4470 17434 4526 17436
rect 4550 17434 4606 17436
rect 4630 17434 4686 17436
rect 4390 17382 4416 17434
rect 4416 17382 4446 17434
rect 4470 17382 4480 17434
rect 4480 17382 4526 17434
rect 4550 17382 4596 17434
rect 4596 17382 4606 17434
rect 4630 17382 4660 17434
rect 4660 17382 4686 17434
rect 4390 17380 4446 17382
rect 4470 17380 4526 17382
rect 4550 17380 4606 17382
rect 4630 17380 4686 17382
rect 7825 17978 7881 17980
rect 7905 17978 7961 17980
rect 7985 17978 8041 17980
rect 8065 17978 8121 17980
rect 7825 17926 7851 17978
rect 7851 17926 7881 17978
rect 7905 17926 7915 17978
rect 7915 17926 7961 17978
rect 7985 17926 8031 17978
rect 8031 17926 8041 17978
rect 8065 17926 8095 17978
rect 8095 17926 8121 17978
rect 7825 17924 7881 17926
rect 7905 17924 7961 17926
rect 7985 17924 8041 17926
rect 8065 17924 8121 17926
rect 7825 16890 7881 16892
rect 7905 16890 7961 16892
rect 7985 16890 8041 16892
rect 8065 16890 8121 16892
rect 7825 16838 7851 16890
rect 7851 16838 7881 16890
rect 7905 16838 7915 16890
rect 7915 16838 7961 16890
rect 7985 16838 8031 16890
rect 8031 16838 8041 16890
rect 8065 16838 8095 16890
rect 8095 16838 8121 16890
rect 7825 16836 7881 16838
rect 7905 16836 7961 16838
rect 7985 16836 8041 16838
rect 8065 16836 8121 16838
rect 4390 16346 4446 16348
rect 4470 16346 4526 16348
rect 4550 16346 4606 16348
rect 4630 16346 4686 16348
rect 4390 16294 4416 16346
rect 4416 16294 4446 16346
rect 4470 16294 4480 16346
rect 4480 16294 4526 16346
rect 4550 16294 4596 16346
rect 4596 16294 4606 16346
rect 4630 16294 4660 16346
rect 4660 16294 4686 16346
rect 4390 16292 4446 16294
rect 4470 16292 4526 16294
rect 4550 16292 4606 16294
rect 4630 16292 4686 16294
rect 7825 15802 7881 15804
rect 7905 15802 7961 15804
rect 7985 15802 8041 15804
rect 8065 15802 8121 15804
rect 7825 15750 7851 15802
rect 7851 15750 7881 15802
rect 7905 15750 7915 15802
rect 7915 15750 7961 15802
rect 7985 15750 8031 15802
rect 8031 15750 8041 15802
rect 8065 15750 8095 15802
rect 8095 15750 8121 15802
rect 7825 15748 7881 15750
rect 7905 15748 7961 15750
rect 7985 15748 8041 15750
rect 8065 15748 8121 15750
rect 4390 15258 4446 15260
rect 4470 15258 4526 15260
rect 4550 15258 4606 15260
rect 4630 15258 4686 15260
rect 4390 15206 4416 15258
rect 4416 15206 4446 15258
rect 4470 15206 4480 15258
rect 4480 15206 4526 15258
rect 4550 15206 4596 15258
rect 4596 15206 4606 15258
rect 4630 15206 4660 15258
rect 4660 15206 4686 15258
rect 4390 15204 4446 15206
rect 4470 15204 4526 15206
rect 4550 15204 4606 15206
rect 4630 15204 4686 15206
rect 7825 14714 7881 14716
rect 7905 14714 7961 14716
rect 7985 14714 8041 14716
rect 8065 14714 8121 14716
rect 7825 14662 7851 14714
rect 7851 14662 7881 14714
rect 7905 14662 7915 14714
rect 7915 14662 7961 14714
rect 7985 14662 8031 14714
rect 8031 14662 8041 14714
rect 8065 14662 8095 14714
rect 8095 14662 8121 14714
rect 7825 14660 7881 14662
rect 7905 14660 7961 14662
rect 7985 14660 8041 14662
rect 8065 14660 8121 14662
rect 4390 14170 4446 14172
rect 4470 14170 4526 14172
rect 4550 14170 4606 14172
rect 4630 14170 4686 14172
rect 4390 14118 4416 14170
rect 4416 14118 4446 14170
rect 4470 14118 4480 14170
rect 4480 14118 4526 14170
rect 4550 14118 4596 14170
rect 4596 14118 4606 14170
rect 4630 14118 4660 14170
rect 4660 14118 4686 14170
rect 4390 14116 4446 14118
rect 4470 14116 4526 14118
rect 4550 14116 4606 14118
rect 4630 14116 4686 14118
rect 3422 13640 3478 13696
rect 7825 13626 7881 13628
rect 7905 13626 7961 13628
rect 7985 13626 8041 13628
rect 8065 13626 8121 13628
rect 7825 13574 7851 13626
rect 7851 13574 7881 13626
rect 7905 13574 7915 13626
rect 7915 13574 7961 13626
rect 7985 13574 8031 13626
rect 8031 13574 8041 13626
rect 8065 13574 8095 13626
rect 8095 13574 8121 13626
rect 7825 13572 7881 13574
rect 7905 13572 7961 13574
rect 7985 13572 8041 13574
rect 8065 13572 8121 13574
rect 4390 13082 4446 13084
rect 4470 13082 4526 13084
rect 4550 13082 4606 13084
rect 4630 13082 4686 13084
rect 4390 13030 4416 13082
rect 4416 13030 4446 13082
rect 4470 13030 4480 13082
rect 4480 13030 4526 13082
rect 4550 13030 4596 13082
rect 4596 13030 4606 13082
rect 4630 13030 4660 13082
rect 4660 13030 4686 13082
rect 4390 13028 4446 13030
rect 4470 13028 4526 13030
rect 4550 13028 4606 13030
rect 4630 13028 4686 13030
rect 7825 12538 7881 12540
rect 7905 12538 7961 12540
rect 7985 12538 8041 12540
rect 8065 12538 8121 12540
rect 7825 12486 7851 12538
rect 7851 12486 7881 12538
rect 7905 12486 7915 12538
rect 7915 12486 7961 12538
rect 7985 12486 8031 12538
rect 8031 12486 8041 12538
rect 8065 12486 8095 12538
rect 8095 12486 8121 12538
rect 7825 12484 7881 12486
rect 7905 12484 7961 12486
rect 7985 12484 8041 12486
rect 8065 12484 8121 12486
rect 4390 11994 4446 11996
rect 4470 11994 4526 11996
rect 4550 11994 4606 11996
rect 4630 11994 4686 11996
rect 4390 11942 4416 11994
rect 4416 11942 4446 11994
rect 4470 11942 4480 11994
rect 4480 11942 4526 11994
rect 4550 11942 4596 11994
rect 4596 11942 4606 11994
rect 4630 11942 4660 11994
rect 4660 11942 4686 11994
rect 4390 11940 4446 11942
rect 4470 11940 4526 11942
rect 4550 11940 4606 11942
rect 4630 11940 4686 11942
rect 7825 11450 7881 11452
rect 7905 11450 7961 11452
rect 7985 11450 8041 11452
rect 8065 11450 8121 11452
rect 7825 11398 7851 11450
rect 7851 11398 7881 11450
rect 7905 11398 7915 11450
rect 7915 11398 7961 11450
rect 7985 11398 8031 11450
rect 8031 11398 8041 11450
rect 8065 11398 8095 11450
rect 8095 11398 8121 11450
rect 7825 11396 7881 11398
rect 7905 11396 7961 11398
rect 7985 11396 8041 11398
rect 8065 11396 8121 11398
rect 4390 10906 4446 10908
rect 4470 10906 4526 10908
rect 4550 10906 4606 10908
rect 4630 10906 4686 10908
rect 4390 10854 4416 10906
rect 4416 10854 4446 10906
rect 4470 10854 4480 10906
rect 4480 10854 4526 10906
rect 4550 10854 4596 10906
rect 4596 10854 4606 10906
rect 4630 10854 4660 10906
rect 4660 10854 4686 10906
rect 4390 10852 4446 10854
rect 4470 10852 4526 10854
rect 4550 10852 4606 10854
rect 4630 10852 4686 10854
rect 7825 10362 7881 10364
rect 7905 10362 7961 10364
rect 7985 10362 8041 10364
rect 8065 10362 8121 10364
rect 7825 10310 7851 10362
rect 7851 10310 7881 10362
rect 7905 10310 7915 10362
rect 7915 10310 7961 10362
rect 7985 10310 8031 10362
rect 8031 10310 8041 10362
rect 8065 10310 8095 10362
rect 8095 10310 8121 10362
rect 7825 10308 7881 10310
rect 7905 10308 7961 10310
rect 7985 10308 8041 10310
rect 8065 10308 8121 10310
rect 4390 9818 4446 9820
rect 4470 9818 4526 9820
rect 4550 9818 4606 9820
rect 4630 9818 4686 9820
rect 4390 9766 4416 9818
rect 4416 9766 4446 9818
rect 4470 9766 4480 9818
rect 4480 9766 4526 9818
rect 4550 9766 4596 9818
rect 4596 9766 4606 9818
rect 4630 9766 4660 9818
rect 4660 9766 4686 9818
rect 4390 9764 4446 9766
rect 4470 9764 4526 9766
rect 4550 9764 4606 9766
rect 4630 9764 4686 9766
rect 4066 9288 4122 9344
rect 7825 9274 7881 9276
rect 7905 9274 7961 9276
rect 7985 9274 8041 9276
rect 8065 9274 8121 9276
rect 7825 9222 7851 9274
rect 7851 9222 7881 9274
rect 7905 9222 7915 9274
rect 7915 9222 7961 9274
rect 7985 9222 8031 9274
rect 8031 9222 8041 9274
rect 8065 9222 8095 9274
rect 8095 9222 8121 9274
rect 7825 9220 7881 9222
rect 7905 9220 7961 9222
rect 7985 9220 8041 9222
rect 8065 9220 8121 9222
rect 11260 21786 11316 21788
rect 11340 21786 11396 21788
rect 11420 21786 11476 21788
rect 11500 21786 11556 21788
rect 11260 21734 11286 21786
rect 11286 21734 11316 21786
rect 11340 21734 11350 21786
rect 11350 21734 11396 21786
rect 11420 21734 11466 21786
rect 11466 21734 11476 21786
rect 11500 21734 11530 21786
rect 11530 21734 11556 21786
rect 11260 21732 11316 21734
rect 11340 21732 11396 21734
rect 11420 21732 11476 21734
rect 11500 21732 11556 21734
rect 14694 22330 14750 22332
rect 14774 22330 14830 22332
rect 14854 22330 14910 22332
rect 14934 22330 14990 22332
rect 14694 22278 14720 22330
rect 14720 22278 14750 22330
rect 14774 22278 14784 22330
rect 14784 22278 14830 22330
rect 14854 22278 14900 22330
rect 14900 22278 14910 22330
rect 14934 22278 14964 22330
rect 14964 22278 14990 22330
rect 14694 22276 14750 22278
rect 14774 22276 14830 22278
rect 14854 22276 14910 22278
rect 14934 22276 14990 22278
rect 11260 20698 11316 20700
rect 11340 20698 11396 20700
rect 11420 20698 11476 20700
rect 11500 20698 11556 20700
rect 11260 20646 11286 20698
rect 11286 20646 11316 20698
rect 11340 20646 11350 20698
rect 11350 20646 11396 20698
rect 11420 20646 11466 20698
rect 11466 20646 11476 20698
rect 11500 20646 11530 20698
rect 11530 20646 11556 20698
rect 11260 20644 11316 20646
rect 11340 20644 11396 20646
rect 11420 20644 11476 20646
rect 11500 20644 11556 20646
rect 11260 19610 11316 19612
rect 11340 19610 11396 19612
rect 11420 19610 11476 19612
rect 11500 19610 11556 19612
rect 11260 19558 11286 19610
rect 11286 19558 11316 19610
rect 11340 19558 11350 19610
rect 11350 19558 11396 19610
rect 11420 19558 11466 19610
rect 11466 19558 11476 19610
rect 11500 19558 11530 19610
rect 11530 19558 11556 19610
rect 11260 19556 11316 19558
rect 11340 19556 11396 19558
rect 11420 19556 11476 19558
rect 11500 19556 11556 19558
rect 11260 18522 11316 18524
rect 11340 18522 11396 18524
rect 11420 18522 11476 18524
rect 11500 18522 11556 18524
rect 11260 18470 11286 18522
rect 11286 18470 11316 18522
rect 11340 18470 11350 18522
rect 11350 18470 11396 18522
rect 11420 18470 11466 18522
rect 11466 18470 11476 18522
rect 11500 18470 11530 18522
rect 11530 18470 11556 18522
rect 11260 18468 11316 18470
rect 11340 18468 11396 18470
rect 11420 18468 11476 18470
rect 11500 18468 11556 18470
rect 11260 17434 11316 17436
rect 11340 17434 11396 17436
rect 11420 17434 11476 17436
rect 11500 17434 11556 17436
rect 11260 17382 11286 17434
rect 11286 17382 11316 17434
rect 11340 17382 11350 17434
rect 11350 17382 11396 17434
rect 11420 17382 11466 17434
rect 11466 17382 11476 17434
rect 11500 17382 11530 17434
rect 11530 17382 11556 17434
rect 11260 17380 11316 17382
rect 11340 17380 11396 17382
rect 11420 17380 11476 17382
rect 11500 17380 11556 17382
rect 11260 16346 11316 16348
rect 11340 16346 11396 16348
rect 11420 16346 11476 16348
rect 11500 16346 11556 16348
rect 11260 16294 11286 16346
rect 11286 16294 11316 16346
rect 11340 16294 11350 16346
rect 11350 16294 11396 16346
rect 11420 16294 11466 16346
rect 11466 16294 11476 16346
rect 11500 16294 11530 16346
rect 11530 16294 11556 16346
rect 11260 16292 11316 16294
rect 11340 16292 11396 16294
rect 11420 16292 11476 16294
rect 11500 16292 11556 16294
rect 11260 15258 11316 15260
rect 11340 15258 11396 15260
rect 11420 15258 11476 15260
rect 11500 15258 11556 15260
rect 11260 15206 11286 15258
rect 11286 15206 11316 15258
rect 11340 15206 11350 15258
rect 11350 15206 11396 15258
rect 11420 15206 11466 15258
rect 11466 15206 11476 15258
rect 11500 15206 11530 15258
rect 11530 15206 11556 15258
rect 11260 15204 11316 15206
rect 11340 15204 11396 15206
rect 11420 15204 11476 15206
rect 11500 15204 11556 15206
rect 11260 14170 11316 14172
rect 11340 14170 11396 14172
rect 11420 14170 11476 14172
rect 11500 14170 11556 14172
rect 11260 14118 11286 14170
rect 11286 14118 11316 14170
rect 11340 14118 11350 14170
rect 11350 14118 11396 14170
rect 11420 14118 11466 14170
rect 11466 14118 11476 14170
rect 11500 14118 11530 14170
rect 11530 14118 11556 14170
rect 11260 14116 11316 14118
rect 11340 14116 11396 14118
rect 11420 14116 11476 14118
rect 11500 14116 11556 14118
rect 11260 13082 11316 13084
rect 11340 13082 11396 13084
rect 11420 13082 11476 13084
rect 11500 13082 11556 13084
rect 11260 13030 11286 13082
rect 11286 13030 11316 13082
rect 11340 13030 11350 13082
rect 11350 13030 11396 13082
rect 11420 13030 11466 13082
rect 11466 13030 11476 13082
rect 11500 13030 11530 13082
rect 11530 13030 11556 13082
rect 11260 13028 11316 13030
rect 11340 13028 11396 13030
rect 11420 13028 11476 13030
rect 11500 13028 11556 13030
rect 11260 11994 11316 11996
rect 11340 11994 11396 11996
rect 11420 11994 11476 11996
rect 11500 11994 11556 11996
rect 11260 11942 11286 11994
rect 11286 11942 11316 11994
rect 11340 11942 11350 11994
rect 11350 11942 11396 11994
rect 11420 11942 11466 11994
rect 11466 11942 11476 11994
rect 11500 11942 11530 11994
rect 11530 11942 11556 11994
rect 11260 11940 11316 11942
rect 11340 11940 11396 11942
rect 11420 11940 11476 11942
rect 11500 11940 11556 11942
rect 11260 10906 11316 10908
rect 11340 10906 11396 10908
rect 11420 10906 11476 10908
rect 11500 10906 11556 10908
rect 11260 10854 11286 10906
rect 11286 10854 11316 10906
rect 11340 10854 11350 10906
rect 11350 10854 11396 10906
rect 11420 10854 11466 10906
rect 11466 10854 11476 10906
rect 11500 10854 11530 10906
rect 11530 10854 11556 10906
rect 11260 10852 11316 10854
rect 11340 10852 11396 10854
rect 11420 10852 11476 10854
rect 11500 10852 11556 10854
rect 11260 9818 11316 9820
rect 11340 9818 11396 9820
rect 11420 9818 11476 9820
rect 11500 9818 11556 9820
rect 11260 9766 11286 9818
rect 11286 9766 11316 9818
rect 11340 9766 11350 9818
rect 11350 9766 11396 9818
rect 11420 9766 11466 9818
rect 11466 9766 11476 9818
rect 11500 9766 11530 9818
rect 11530 9766 11556 9818
rect 11260 9764 11316 9766
rect 11340 9764 11396 9766
rect 11420 9764 11476 9766
rect 11500 9764 11556 9766
rect 4390 8730 4446 8732
rect 4470 8730 4526 8732
rect 4550 8730 4606 8732
rect 4630 8730 4686 8732
rect 4390 8678 4416 8730
rect 4416 8678 4446 8730
rect 4470 8678 4480 8730
rect 4480 8678 4526 8730
rect 4550 8678 4596 8730
rect 4596 8678 4606 8730
rect 4630 8678 4660 8730
rect 4660 8678 4686 8730
rect 4390 8676 4446 8678
rect 4470 8676 4526 8678
rect 4550 8676 4606 8678
rect 4630 8676 4686 8678
rect 11260 8730 11316 8732
rect 11340 8730 11396 8732
rect 11420 8730 11476 8732
rect 11500 8730 11556 8732
rect 11260 8678 11286 8730
rect 11286 8678 11316 8730
rect 11340 8678 11350 8730
rect 11350 8678 11396 8730
rect 11420 8678 11466 8730
rect 11466 8678 11476 8730
rect 11500 8678 11530 8730
rect 11530 8678 11556 8730
rect 11260 8676 11316 8678
rect 11340 8676 11396 8678
rect 11420 8676 11476 8678
rect 11500 8676 11556 8678
rect 7825 8186 7881 8188
rect 7905 8186 7961 8188
rect 7985 8186 8041 8188
rect 8065 8186 8121 8188
rect 7825 8134 7851 8186
rect 7851 8134 7881 8186
rect 7905 8134 7915 8186
rect 7915 8134 7961 8186
rect 7985 8134 8031 8186
rect 8031 8134 8041 8186
rect 8065 8134 8095 8186
rect 8095 8134 8121 8186
rect 7825 8132 7881 8134
rect 7905 8132 7961 8134
rect 7985 8132 8041 8134
rect 8065 8132 8121 8134
rect 4390 7642 4446 7644
rect 4470 7642 4526 7644
rect 4550 7642 4606 7644
rect 4630 7642 4686 7644
rect 4390 7590 4416 7642
rect 4416 7590 4446 7642
rect 4470 7590 4480 7642
rect 4480 7590 4526 7642
rect 4550 7590 4596 7642
rect 4596 7590 4606 7642
rect 4630 7590 4660 7642
rect 4660 7590 4686 7642
rect 4390 7588 4446 7590
rect 4470 7588 4526 7590
rect 4550 7588 4606 7590
rect 4630 7588 4686 7590
rect 11260 7642 11316 7644
rect 11340 7642 11396 7644
rect 11420 7642 11476 7644
rect 11500 7642 11556 7644
rect 11260 7590 11286 7642
rect 11286 7590 11316 7642
rect 11340 7590 11350 7642
rect 11350 7590 11396 7642
rect 11420 7590 11466 7642
rect 11466 7590 11476 7642
rect 11500 7590 11530 7642
rect 11530 7590 11556 7642
rect 11260 7588 11316 7590
rect 11340 7588 11396 7590
rect 11420 7588 11476 7590
rect 11500 7588 11556 7590
rect 7825 7098 7881 7100
rect 7905 7098 7961 7100
rect 7985 7098 8041 7100
rect 8065 7098 8121 7100
rect 7825 7046 7851 7098
rect 7851 7046 7881 7098
rect 7905 7046 7915 7098
rect 7915 7046 7961 7098
rect 7985 7046 8031 7098
rect 8031 7046 8041 7098
rect 8065 7046 8095 7098
rect 8095 7046 8121 7098
rect 7825 7044 7881 7046
rect 7905 7044 7961 7046
rect 7985 7044 8041 7046
rect 8065 7044 8121 7046
rect 4390 6554 4446 6556
rect 4470 6554 4526 6556
rect 4550 6554 4606 6556
rect 4630 6554 4686 6556
rect 4390 6502 4416 6554
rect 4416 6502 4446 6554
rect 4470 6502 4480 6554
rect 4480 6502 4526 6554
rect 4550 6502 4596 6554
rect 4596 6502 4606 6554
rect 4630 6502 4660 6554
rect 4660 6502 4686 6554
rect 4390 6500 4446 6502
rect 4470 6500 4526 6502
rect 4550 6500 4606 6502
rect 4630 6500 4686 6502
rect 11260 6554 11316 6556
rect 11340 6554 11396 6556
rect 11420 6554 11476 6556
rect 11500 6554 11556 6556
rect 11260 6502 11286 6554
rect 11286 6502 11316 6554
rect 11340 6502 11350 6554
rect 11350 6502 11396 6554
rect 11420 6502 11466 6554
rect 11466 6502 11476 6554
rect 11500 6502 11530 6554
rect 11530 6502 11556 6554
rect 11260 6500 11316 6502
rect 11340 6500 11396 6502
rect 11420 6500 11476 6502
rect 11500 6500 11556 6502
rect 7825 6010 7881 6012
rect 7905 6010 7961 6012
rect 7985 6010 8041 6012
rect 8065 6010 8121 6012
rect 7825 5958 7851 6010
rect 7851 5958 7881 6010
rect 7905 5958 7915 6010
rect 7915 5958 7961 6010
rect 7985 5958 8031 6010
rect 8031 5958 8041 6010
rect 8065 5958 8095 6010
rect 8095 5958 8121 6010
rect 7825 5956 7881 5958
rect 7905 5956 7961 5958
rect 7985 5956 8041 5958
rect 8065 5956 8121 5958
rect 4390 5466 4446 5468
rect 4470 5466 4526 5468
rect 4550 5466 4606 5468
rect 4630 5466 4686 5468
rect 4390 5414 4416 5466
rect 4416 5414 4446 5466
rect 4470 5414 4480 5466
rect 4480 5414 4526 5466
rect 4550 5414 4596 5466
rect 4596 5414 4606 5466
rect 4630 5414 4660 5466
rect 4660 5414 4686 5466
rect 4390 5412 4446 5414
rect 4470 5412 4526 5414
rect 4550 5412 4606 5414
rect 4630 5412 4686 5414
rect 11260 5466 11316 5468
rect 11340 5466 11396 5468
rect 11420 5466 11476 5468
rect 11500 5466 11556 5468
rect 11260 5414 11286 5466
rect 11286 5414 11316 5466
rect 11340 5414 11350 5466
rect 11350 5414 11396 5466
rect 11420 5414 11466 5466
rect 11466 5414 11476 5466
rect 11500 5414 11530 5466
rect 11530 5414 11556 5466
rect 11260 5412 11316 5414
rect 11340 5412 11396 5414
rect 11420 5412 11476 5414
rect 11500 5412 11556 5414
rect 7825 4922 7881 4924
rect 7905 4922 7961 4924
rect 7985 4922 8041 4924
rect 8065 4922 8121 4924
rect 7825 4870 7851 4922
rect 7851 4870 7881 4922
rect 7905 4870 7915 4922
rect 7915 4870 7961 4922
rect 7985 4870 8031 4922
rect 8031 4870 8041 4922
rect 8065 4870 8095 4922
rect 8095 4870 8121 4922
rect 7825 4868 7881 4870
rect 7905 4868 7961 4870
rect 7985 4868 8041 4870
rect 8065 4868 8121 4870
rect 4390 4378 4446 4380
rect 4470 4378 4526 4380
rect 4550 4378 4606 4380
rect 4630 4378 4686 4380
rect 4390 4326 4416 4378
rect 4416 4326 4446 4378
rect 4470 4326 4480 4378
rect 4480 4326 4526 4378
rect 4550 4326 4596 4378
rect 4596 4326 4606 4378
rect 4630 4326 4660 4378
rect 4660 4326 4686 4378
rect 4390 4324 4446 4326
rect 4470 4324 4526 4326
rect 4550 4324 4606 4326
rect 4630 4324 4686 4326
rect 11260 4378 11316 4380
rect 11340 4378 11396 4380
rect 11420 4378 11476 4380
rect 11500 4378 11556 4380
rect 11260 4326 11286 4378
rect 11286 4326 11316 4378
rect 11340 4326 11350 4378
rect 11350 4326 11396 4378
rect 11420 4326 11466 4378
rect 11466 4326 11476 4378
rect 11500 4326 11530 4378
rect 11530 4326 11556 4378
rect 11260 4324 11316 4326
rect 11340 4324 11396 4326
rect 11420 4324 11476 4326
rect 11500 4324 11556 4326
rect 4390 3290 4446 3292
rect 4470 3290 4526 3292
rect 4550 3290 4606 3292
rect 4630 3290 4686 3292
rect 4390 3238 4416 3290
rect 4416 3238 4446 3290
rect 4470 3238 4480 3290
rect 4480 3238 4526 3290
rect 4550 3238 4596 3290
rect 4596 3238 4606 3290
rect 4630 3238 4660 3290
rect 4660 3238 4686 3290
rect 4390 3236 4446 3238
rect 4470 3236 4526 3238
rect 4550 3236 4606 3238
rect 4630 3236 4686 3238
rect 4390 2202 4446 2204
rect 4470 2202 4526 2204
rect 4550 2202 4606 2204
rect 4630 2202 4686 2204
rect 4390 2150 4416 2202
rect 4416 2150 4446 2202
rect 4470 2150 4480 2202
rect 4480 2150 4526 2202
rect 4550 2150 4596 2202
rect 4596 2150 4606 2202
rect 4630 2150 4660 2202
rect 4660 2150 4686 2202
rect 4390 2148 4446 2150
rect 4470 2148 4526 2150
rect 4550 2148 4606 2150
rect 4630 2148 4686 2150
rect 7825 3834 7881 3836
rect 7905 3834 7961 3836
rect 7985 3834 8041 3836
rect 8065 3834 8121 3836
rect 7825 3782 7851 3834
rect 7851 3782 7881 3834
rect 7905 3782 7915 3834
rect 7915 3782 7961 3834
rect 7985 3782 8031 3834
rect 8031 3782 8041 3834
rect 8065 3782 8095 3834
rect 8095 3782 8121 3834
rect 7825 3780 7881 3782
rect 7905 3780 7961 3782
rect 7985 3780 8041 3782
rect 8065 3780 8121 3782
rect 7825 2746 7881 2748
rect 7905 2746 7961 2748
rect 7985 2746 8041 2748
rect 8065 2746 8121 2748
rect 7825 2694 7851 2746
rect 7851 2694 7881 2746
rect 7905 2694 7915 2746
rect 7915 2694 7961 2746
rect 7985 2694 8031 2746
rect 8031 2694 8041 2746
rect 8065 2694 8095 2746
rect 8095 2694 8121 2746
rect 7825 2692 7881 2694
rect 7905 2692 7961 2694
rect 7985 2692 8041 2694
rect 8065 2692 8121 2694
rect 14694 21242 14750 21244
rect 14774 21242 14830 21244
rect 14854 21242 14910 21244
rect 14934 21242 14990 21244
rect 14694 21190 14720 21242
rect 14720 21190 14750 21242
rect 14774 21190 14784 21242
rect 14784 21190 14830 21242
rect 14854 21190 14900 21242
rect 14900 21190 14910 21242
rect 14934 21190 14964 21242
rect 14964 21190 14990 21242
rect 14694 21188 14750 21190
rect 14774 21188 14830 21190
rect 14854 21188 14910 21190
rect 14934 21188 14990 21190
rect 14694 20154 14750 20156
rect 14774 20154 14830 20156
rect 14854 20154 14910 20156
rect 14934 20154 14990 20156
rect 14694 20102 14720 20154
rect 14720 20102 14750 20154
rect 14774 20102 14784 20154
rect 14784 20102 14830 20154
rect 14854 20102 14900 20154
rect 14900 20102 14910 20154
rect 14934 20102 14964 20154
rect 14964 20102 14990 20154
rect 14694 20100 14750 20102
rect 14774 20100 14830 20102
rect 14854 20100 14910 20102
rect 14934 20100 14990 20102
rect 14694 19066 14750 19068
rect 14774 19066 14830 19068
rect 14854 19066 14910 19068
rect 14934 19066 14990 19068
rect 14694 19014 14720 19066
rect 14720 19014 14750 19066
rect 14774 19014 14784 19066
rect 14784 19014 14830 19066
rect 14854 19014 14900 19066
rect 14900 19014 14910 19066
rect 14934 19014 14964 19066
rect 14964 19014 14990 19066
rect 14694 19012 14750 19014
rect 14774 19012 14830 19014
rect 14854 19012 14910 19014
rect 14934 19012 14990 19014
rect 14694 17978 14750 17980
rect 14774 17978 14830 17980
rect 14854 17978 14910 17980
rect 14934 17978 14990 17980
rect 14694 17926 14720 17978
rect 14720 17926 14750 17978
rect 14774 17926 14784 17978
rect 14784 17926 14830 17978
rect 14854 17926 14900 17978
rect 14900 17926 14910 17978
rect 14934 17926 14964 17978
rect 14964 17926 14990 17978
rect 14694 17924 14750 17926
rect 14774 17924 14830 17926
rect 14854 17924 14910 17926
rect 14934 17924 14990 17926
rect 14694 16890 14750 16892
rect 14774 16890 14830 16892
rect 14854 16890 14910 16892
rect 14934 16890 14990 16892
rect 14694 16838 14720 16890
rect 14720 16838 14750 16890
rect 14774 16838 14784 16890
rect 14784 16838 14830 16890
rect 14854 16838 14900 16890
rect 14900 16838 14910 16890
rect 14934 16838 14964 16890
rect 14964 16838 14990 16890
rect 14694 16836 14750 16838
rect 14774 16836 14830 16838
rect 14854 16836 14910 16838
rect 14934 16836 14990 16838
rect 14694 15802 14750 15804
rect 14774 15802 14830 15804
rect 14854 15802 14910 15804
rect 14934 15802 14990 15804
rect 14694 15750 14720 15802
rect 14720 15750 14750 15802
rect 14774 15750 14784 15802
rect 14784 15750 14830 15802
rect 14854 15750 14900 15802
rect 14900 15750 14910 15802
rect 14934 15750 14964 15802
rect 14964 15750 14990 15802
rect 14694 15748 14750 15750
rect 14774 15748 14830 15750
rect 14854 15748 14910 15750
rect 14934 15748 14990 15750
rect 14694 14714 14750 14716
rect 14774 14714 14830 14716
rect 14854 14714 14910 14716
rect 14934 14714 14990 14716
rect 14694 14662 14720 14714
rect 14720 14662 14750 14714
rect 14774 14662 14784 14714
rect 14784 14662 14830 14714
rect 14854 14662 14900 14714
rect 14900 14662 14910 14714
rect 14934 14662 14964 14714
rect 14964 14662 14990 14714
rect 14694 14660 14750 14662
rect 14774 14660 14830 14662
rect 14854 14660 14910 14662
rect 14934 14660 14990 14662
rect 14694 13626 14750 13628
rect 14774 13626 14830 13628
rect 14854 13626 14910 13628
rect 14934 13626 14990 13628
rect 14694 13574 14720 13626
rect 14720 13574 14750 13626
rect 14774 13574 14784 13626
rect 14784 13574 14830 13626
rect 14854 13574 14900 13626
rect 14900 13574 14910 13626
rect 14934 13574 14964 13626
rect 14964 13574 14990 13626
rect 14694 13572 14750 13574
rect 14774 13572 14830 13574
rect 14854 13572 14910 13574
rect 14934 13572 14990 13574
rect 14694 12538 14750 12540
rect 14774 12538 14830 12540
rect 14854 12538 14910 12540
rect 14934 12538 14990 12540
rect 14694 12486 14720 12538
rect 14720 12486 14750 12538
rect 14774 12486 14784 12538
rect 14784 12486 14830 12538
rect 14854 12486 14900 12538
rect 14900 12486 14910 12538
rect 14934 12486 14964 12538
rect 14964 12486 14990 12538
rect 14694 12484 14750 12486
rect 14774 12484 14830 12486
rect 14854 12484 14910 12486
rect 14934 12484 14990 12486
rect 14694 11450 14750 11452
rect 14774 11450 14830 11452
rect 14854 11450 14910 11452
rect 14934 11450 14990 11452
rect 14694 11398 14720 11450
rect 14720 11398 14750 11450
rect 14774 11398 14784 11450
rect 14784 11398 14830 11450
rect 14854 11398 14900 11450
rect 14900 11398 14910 11450
rect 14934 11398 14964 11450
rect 14964 11398 14990 11450
rect 14694 11396 14750 11398
rect 14774 11396 14830 11398
rect 14854 11396 14910 11398
rect 14934 11396 14990 11398
rect 18129 21786 18185 21788
rect 18209 21786 18265 21788
rect 18289 21786 18345 21788
rect 18369 21786 18425 21788
rect 18129 21734 18155 21786
rect 18155 21734 18185 21786
rect 18209 21734 18219 21786
rect 18219 21734 18265 21786
rect 18289 21734 18335 21786
rect 18335 21734 18345 21786
rect 18369 21734 18399 21786
rect 18399 21734 18425 21786
rect 18129 21732 18185 21734
rect 18209 21732 18265 21734
rect 18289 21732 18345 21734
rect 18369 21732 18425 21734
rect 18129 20698 18185 20700
rect 18209 20698 18265 20700
rect 18289 20698 18345 20700
rect 18369 20698 18425 20700
rect 18129 20646 18155 20698
rect 18155 20646 18185 20698
rect 18209 20646 18219 20698
rect 18219 20646 18265 20698
rect 18289 20646 18335 20698
rect 18335 20646 18345 20698
rect 18369 20646 18399 20698
rect 18399 20646 18425 20698
rect 18129 20644 18185 20646
rect 18209 20644 18265 20646
rect 18289 20644 18345 20646
rect 18369 20644 18425 20646
rect 18418 19896 18474 19952
rect 18129 19610 18185 19612
rect 18209 19610 18265 19612
rect 18289 19610 18345 19612
rect 18369 19610 18425 19612
rect 18129 19558 18155 19610
rect 18155 19558 18185 19610
rect 18209 19558 18219 19610
rect 18219 19558 18265 19610
rect 18289 19558 18335 19610
rect 18335 19558 18345 19610
rect 18369 19558 18399 19610
rect 18399 19558 18425 19610
rect 18129 19556 18185 19558
rect 18209 19556 18265 19558
rect 18289 19556 18345 19558
rect 18369 19556 18425 19558
rect 18129 18522 18185 18524
rect 18209 18522 18265 18524
rect 18289 18522 18345 18524
rect 18369 18522 18425 18524
rect 18129 18470 18155 18522
rect 18155 18470 18185 18522
rect 18209 18470 18219 18522
rect 18219 18470 18265 18522
rect 18289 18470 18335 18522
rect 18335 18470 18345 18522
rect 18369 18470 18399 18522
rect 18399 18470 18425 18522
rect 18129 18468 18185 18470
rect 18209 18468 18265 18470
rect 18289 18468 18345 18470
rect 18369 18468 18425 18470
rect 18129 17434 18185 17436
rect 18209 17434 18265 17436
rect 18289 17434 18345 17436
rect 18369 17434 18425 17436
rect 18129 17382 18155 17434
rect 18155 17382 18185 17434
rect 18209 17382 18219 17434
rect 18219 17382 18265 17434
rect 18289 17382 18335 17434
rect 18335 17382 18345 17434
rect 18369 17382 18399 17434
rect 18399 17382 18425 17434
rect 18129 17380 18185 17382
rect 18209 17380 18265 17382
rect 18289 17380 18345 17382
rect 18369 17380 18425 17382
rect 18129 16346 18185 16348
rect 18209 16346 18265 16348
rect 18289 16346 18345 16348
rect 18369 16346 18425 16348
rect 18129 16294 18155 16346
rect 18155 16294 18185 16346
rect 18209 16294 18219 16346
rect 18219 16294 18265 16346
rect 18289 16294 18335 16346
rect 18335 16294 18345 16346
rect 18369 16294 18399 16346
rect 18399 16294 18425 16346
rect 18129 16292 18185 16294
rect 18209 16292 18265 16294
rect 18289 16292 18345 16294
rect 18369 16292 18425 16294
rect 19522 15544 19578 15600
rect 18129 15258 18185 15260
rect 18209 15258 18265 15260
rect 18289 15258 18345 15260
rect 18369 15258 18425 15260
rect 18129 15206 18155 15258
rect 18155 15206 18185 15258
rect 18209 15206 18219 15258
rect 18219 15206 18265 15258
rect 18289 15206 18335 15258
rect 18335 15206 18345 15258
rect 18369 15206 18399 15258
rect 18399 15206 18425 15258
rect 18129 15204 18185 15206
rect 18209 15204 18265 15206
rect 18289 15204 18345 15206
rect 18369 15204 18425 15206
rect 18129 14170 18185 14172
rect 18209 14170 18265 14172
rect 18289 14170 18345 14172
rect 18369 14170 18425 14172
rect 18129 14118 18155 14170
rect 18155 14118 18185 14170
rect 18209 14118 18219 14170
rect 18219 14118 18265 14170
rect 18289 14118 18335 14170
rect 18335 14118 18345 14170
rect 18369 14118 18399 14170
rect 18399 14118 18425 14170
rect 18129 14116 18185 14118
rect 18209 14116 18265 14118
rect 18289 14116 18345 14118
rect 18369 14116 18425 14118
rect 18129 13082 18185 13084
rect 18209 13082 18265 13084
rect 18289 13082 18345 13084
rect 18369 13082 18425 13084
rect 18129 13030 18155 13082
rect 18155 13030 18185 13082
rect 18209 13030 18219 13082
rect 18219 13030 18265 13082
rect 18289 13030 18335 13082
rect 18335 13030 18345 13082
rect 18369 13030 18399 13082
rect 18399 13030 18425 13082
rect 18129 13028 18185 13030
rect 18209 13028 18265 13030
rect 18289 13028 18345 13030
rect 18369 13028 18425 13030
rect 14694 10362 14750 10364
rect 14774 10362 14830 10364
rect 14854 10362 14910 10364
rect 14934 10362 14990 10364
rect 14694 10310 14720 10362
rect 14720 10310 14750 10362
rect 14774 10310 14784 10362
rect 14784 10310 14830 10362
rect 14854 10310 14900 10362
rect 14900 10310 14910 10362
rect 14934 10310 14964 10362
rect 14964 10310 14990 10362
rect 14694 10308 14750 10310
rect 14774 10308 14830 10310
rect 14854 10308 14910 10310
rect 14934 10308 14990 10310
rect 14694 9274 14750 9276
rect 14774 9274 14830 9276
rect 14854 9274 14910 9276
rect 14934 9274 14990 9276
rect 14694 9222 14720 9274
rect 14720 9222 14750 9274
rect 14774 9222 14784 9274
rect 14784 9222 14830 9274
rect 14854 9222 14900 9274
rect 14900 9222 14910 9274
rect 14934 9222 14964 9274
rect 14964 9222 14990 9274
rect 14694 9220 14750 9222
rect 14774 9220 14830 9222
rect 14854 9220 14910 9222
rect 14934 9220 14990 9222
rect 11260 3290 11316 3292
rect 11340 3290 11396 3292
rect 11420 3290 11476 3292
rect 11500 3290 11556 3292
rect 11260 3238 11286 3290
rect 11286 3238 11316 3290
rect 11340 3238 11350 3290
rect 11350 3238 11396 3290
rect 11420 3238 11466 3290
rect 11466 3238 11476 3290
rect 11500 3238 11530 3290
rect 11530 3238 11556 3290
rect 11260 3236 11316 3238
rect 11340 3236 11396 3238
rect 11420 3236 11476 3238
rect 11500 3236 11556 3238
rect 11260 2202 11316 2204
rect 11340 2202 11396 2204
rect 11420 2202 11476 2204
rect 11500 2202 11556 2204
rect 11260 2150 11286 2202
rect 11286 2150 11316 2202
rect 11340 2150 11350 2202
rect 11350 2150 11396 2202
rect 11420 2150 11466 2202
rect 11466 2150 11476 2202
rect 11500 2150 11530 2202
rect 11530 2150 11556 2202
rect 11260 2148 11316 2150
rect 11340 2148 11396 2150
rect 11420 2148 11476 2150
rect 11500 2148 11556 2150
rect 14694 8186 14750 8188
rect 14774 8186 14830 8188
rect 14854 8186 14910 8188
rect 14934 8186 14990 8188
rect 14694 8134 14720 8186
rect 14720 8134 14750 8186
rect 14774 8134 14784 8186
rect 14784 8134 14830 8186
rect 14854 8134 14900 8186
rect 14900 8134 14910 8186
rect 14934 8134 14964 8186
rect 14964 8134 14990 8186
rect 14694 8132 14750 8134
rect 14774 8132 14830 8134
rect 14854 8132 14910 8134
rect 14934 8132 14990 8134
rect 14694 7098 14750 7100
rect 14774 7098 14830 7100
rect 14854 7098 14910 7100
rect 14934 7098 14990 7100
rect 14694 7046 14720 7098
rect 14720 7046 14750 7098
rect 14774 7046 14784 7098
rect 14784 7046 14830 7098
rect 14854 7046 14900 7098
rect 14900 7046 14910 7098
rect 14934 7046 14964 7098
rect 14964 7046 14990 7098
rect 14694 7044 14750 7046
rect 14774 7044 14830 7046
rect 14854 7044 14910 7046
rect 14934 7044 14990 7046
rect 14694 6010 14750 6012
rect 14774 6010 14830 6012
rect 14854 6010 14910 6012
rect 14934 6010 14990 6012
rect 14694 5958 14720 6010
rect 14720 5958 14750 6010
rect 14774 5958 14784 6010
rect 14784 5958 14830 6010
rect 14854 5958 14900 6010
rect 14900 5958 14910 6010
rect 14934 5958 14964 6010
rect 14964 5958 14990 6010
rect 14694 5956 14750 5958
rect 14774 5956 14830 5958
rect 14854 5956 14910 5958
rect 14934 5956 14990 5958
rect 14694 4922 14750 4924
rect 14774 4922 14830 4924
rect 14854 4922 14910 4924
rect 14934 4922 14990 4924
rect 14694 4870 14720 4922
rect 14720 4870 14750 4922
rect 14774 4870 14784 4922
rect 14784 4870 14830 4922
rect 14854 4870 14900 4922
rect 14900 4870 14910 4922
rect 14934 4870 14964 4922
rect 14964 4870 14990 4922
rect 14694 4868 14750 4870
rect 14774 4868 14830 4870
rect 14854 4868 14910 4870
rect 14934 4868 14990 4870
rect 14694 3834 14750 3836
rect 14774 3834 14830 3836
rect 14854 3834 14910 3836
rect 14934 3834 14990 3836
rect 14694 3782 14720 3834
rect 14720 3782 14750 3834
rect 14774 3782 14784 3834
rect 14784 3782 14830 3834
rect 14854 3782 14900 3834
rect 14900 3782 14910 3834
rect 14934 3782 14964 3834
rect 14964 3782 14990 3834
rect 14694 3780 14750 3782
rect 14774 3780 14830 3782
rect 14854 3780 14910 3782
rect 14934 3780 14990 3782
rect 14694 2746 14750 2748
rect 14774 2746 14830 2748
rect 14854 2746 14910 2748
rect 14934 2746 14990 2748
rect 14694 2694 14720 2746
rect 14720 2694 14750 2746
rect 14774 2694 14784 2746
rect 14784 2694 14830 2746
rect 14854 2694 14900 2746
rect 14900 2694 14910 2746
rect 14934 2694 14964 2746
rect 14964 2694 14990 2746
rect 14694 2692 14750 2694
rect 14774 2692 14830 2694
rect 14854 2692 14910 2694
rect 14934 2692 14990 2694
rect 18129 11994 18185 11996
rect 18209 11994 18265 11996
rect 18289 11994 18345 11996
rect 18369 11994 18425 11996
rect 18129 11942 18155 11994
rect 18155 11942 18185 11994
rect 18209 11942 18219 11994
rect 18219 11942 18265 11994
rect 18289 11942 18335 11994
rect 18335 11942 18345 11994
rect 18369 11942 18399 11994
rect 18399 11942 18425 11994
rect 18129 11940 18185 11942
rect 18209 11940 18265 11942
rect 18289 11940 18345 11942
rect 18369 11940 18425 11942
rect 18129 10906 18185 10908
rect 18209 10906 18265 10908
rect 18289 10906 18345 10908
rect 18369 10906 18425 10908
rect 18129 10854 18155 10906
rect 18155 10854 18185 10906
rect 18209 10854 18219 10906
rect 18219 10854 18265 10906
rect 18289 10854 18335 10906
rect 18335 10854 18345 10906
rect 18369 10854 18399 10906
rect 18399 10854 18425 10906
rect 18129 10852 18185 10854
rect 18209 10852 18265 10854
rect 18289 10852 18345 10854
rect 18369 10852 18425 10854
rect 19706 11192 19762 11248
rect 18129 9818 18185 9820
rect 18209 9818 18265 9820
rect 18289 9818 18345 9820
rect 18369 9818 18425 9820
rect 18129 9766 18155 9818
rect 18155 9766 18185 9818
rect 18209 9766 18219 9818
rect 18219 9766 18265 9818
rect 18289 9766 18335 9818
rect 18335 9766 18345 9818
rect 18369 9766 18399 9818
rect 18399 9766 18425 9818
rect 18129 9764 18185 9766
rect 18209 9764 18265 9766
rect 18289 9764 18345 9766
rect 18369 9764 18425 9766
rect 18129 8730 18185 8732
rect 18209 8730 18265 8732
rect 18289 8730 18345 8732
rect 18369 8730 18425 8732
rect 18129 8678 18155 8730
rect 18155 8678 18185 8730
rect 18209 8678 18219 8730
rect 18219 8678 18265 8730
rect 18289 8678 18335 8730
rect 18335 8678 18345 8730
rect 18369 8678 18399 8730
rect 18399 8678 18425 8730
rect 18129 8676 18185 8678
rect 18209 8676 18265 8678
rect 18289 8676 18345 8678
rect 18369 8676 18425 8678
rect 18129 7642 18185 7644
rect 18209 7642 18265 7644
rect 18289 7642 18345 7644
rect 18369 7642 18425 7644
rect 18129 7590 18155 7642
rect 18155 7590 18185 7642
rect 18209 7590 18219 7642
rect 18219 7590 18265 7642
rect 18289 7590 18335 7642
rect 18335 7590 18345 7642
rect 18369 7590 18399 7642
rect 18399 7590 18425 7642
rect 18129 7588 18185 7590
rect 18209 7588 18265 7590
rect 18289 7588 18345 7590
rect 18369 7588 18425 7590
rect 19982 7112 20038 7168
rect 18129 6554 18185 6556
rect 18209 6554 18265 6556
rect 18289 6554 18345 6556
rect 18369 6554 18425 6556
rect 18129 6502 18155 6554
rect 18155 6502 18185 6554
rect 18209 6502 18219 6554
rect 18219 6502 18265 6554
rect 18289 6502 18335 6554
rect 18335 6502 18345 6554
rect 18369 6502 18399 6554
rect 18399 6502 18425 6554
rect 18129 6500 18185 6502
rect 18209 6500 18265 6502
rect 18289 6500 18345 6502
rect 18369 6500 18425 6502
rect 18129 5466 18185 5468
rect 18209 5466 18265 5468
rect 18289 5466 18345 5468
rect 18369 5466 18425 5468
rect 18129 5414 18155 5466
rect 18155 5414 18185 5466
rect 18209 5414 18219 5466
rect 18219 5414 18265 5466
rect 18289 5414 18335 5466
rect 18335 5414 18345 5466
rect 18369 5414 18399 5466
rect 18399 5414 18425 5466
rect 18129 5412 18185 5414
rect 18209 5412 18265 5414
rect 18289 5412 18345 5414
rect 18369 5412 18425 5414
rect 18129 4378 18185 4380
rect 18209 4378 18265 4380
rect 18289 4378 18345 4380
rect 18369 4378 18425 4380
rect 18129 4326 18155 4378
rect 18155 4326 18185 4378
rect 18209 4326 18219 4378
rect 18219 4326 18265 4378
rect 18289 4326 18335 4378
rect 18335 4326 18345 4378
rect 18369 4326 18399 4378
rect 18399 4326 18425 4378
rect 18129 4324 18185 4326
rect 18209 4324 18265 4326
rect 18289 4324 18345 4326
rect 18369 4324 18425 4326
rect 18129 3290 18185 3292
rect 18209 3290 18265 3292
rect 18289 3290 18345 3292
rect 18369 3290 18425 3292
rect 18129 3238 18155 3290
rect 18155 3238 18185 3290
rect 18209 3238 18219 3290
rect 18219 3238 18265 3290
rect 18289 3238 18335 3290
rect 18335 3238 18345 3290
rect 18369 3238 18399 3290
rect 18399 3238 18425 3290
rect 18129 3236 18185 3238
rect 18209 3236 18265 3238
rect 18289 3236 18345 3238
rect 18369 3236 18425 3238
rect 20350 2760 20406 2816
rect 18129 2202 18185 2204
rect 18209 2202 18265 2204
rect 18289 2202 18345 2204
rect 18369 2202 18425 2204
rect 18129 2150 18155 2202
rect 18155 2150 18185 2202
rect 18209 2150 18219 2202
rect 18219 2150 18265 2202
rect 18289 2150 18335 2202
rect 18335 2150 18345 2202
rect 18369 2150 18399 2202
rect 18399 2150 18425 2202
rect 18129 2148 18185 2150
rect 18209 2148 18265 2150
rect 18289 2148 18345 2150
rect 18369 2148 18425 2150
<< metal3 >>
rect 7813 22336 8133 22337
rect 7813 22272 7821 22336
rect 7885 22272 7901 22336
rect 7965 22272 7981 22336
rect 8045 22272 8061 22336
rect 8125 22272 8133 22336
rect 7813 22271 8133 22272
rect 14682 22336 15002 22337
rect 14682 22272 14690 22336
rect 14754 22272 14770 22336
rect 14834 22272 14850 22336
rect 14914 22272 14930 22336
rect 14994 22272 15002 22336
rect 14682 22271 15002 22272
rect 0 22130 800 22160
rect 1577 22130 1643 22133
rect 0 22128 1643 22130
rect 0 22072 1582 22128
rect 1638 22072 1643 22128
rect 0 22070 1643 22072
rect 0 22040 800 22070
rect 1577 22067 1643 22070
rect 4378 21792 4698 21793
rect 4378 21728 4386 21792
rect 4450 21728 4466 21792
rect 4530 21728 4546 21792
rect 4610 21728 4626 21792
rect 4690 21728 4698 21792
rect 4378 21727 4698 21728
rect 11248 21792 11568 21793
rect 11248 21728 11256 21792
rect 11320 21728 11336 21792
rect 11400 21728 11416 21792
rect 11480 21728 11496 21792
rect 11560 21728 11568 21792
rect 11248 21727 11568 21728
rect 18117 21792 18437 21793
rect 18117 21728 18125 21792
rect 18189 21728 18205 21792
rect 18269 21728 18285 21792
rect 18349 21728 18365 21792
rect 18429 21728 18437 21792
rect 18117 21727 18437 21728
rect 7813 21248 8133 21249
rect 7813 21184 7821 21248
rect 7885 21184 7901 21248
rect 7965 21184 7981 21248
rect 8045 21184 8061 21248
rect 8125 21184 8133 21248
rect 7813 21183 8133 21184
rect 14682 21248 15002 21249
rect 14682 21184 14690 21248
rect 14754 21184 14770 21248
rect 14834 21184 14850 21248
rect 14914 21184 14930 21248
rect 14994 21184 15002 21248
rect 14682 21183 15002 21184
rect 4378 20704 4698 20705
rect 4378 20640 4386 20704
rect 4450 20640 4466 20704
rect 4530 20640 4546 20704
rect 4610 20640 4626 20704
rect 4690 20640 4698 20704
rect 4378 20639 4698 20640
rect 11248 20704 11568 20705
rect 11248 20640 11256 20704
rect 11320 20640 11336 20704
rect 11400 20640 11416 20704
rect 11480 20640 11496 20704
rect 11560 20640 11568 20704
rect 11248 20639 11568 20640
rect 18117 20704 18437 20705
rect 18117 20640 18125 20704
rect 18189 20640 18205 20704
rect 18269 20640 18285 20704
rect 18349 20640 18365 20704
rect 18429 20640 18437 20704
rect 18117 20639 18437 20640
rect 7813 20160 8133 20161
rect 7813 20096 7821 20160
rect 7885 20096 7901 20160
rect 7965 20096 7981 20160
rect 8045 20096 8061 20160
rect 8125 20096 8133 20160
rect 7813 20095 8133 20096
rect 14682 20160 15002 20161
rect 14682 20096 14690 20160
rect 14754 20096 14770 20160
rect 14834 20096 14850 20160
rect 14914 20096 14930 20160
rect 14994 20096 15002 20160
rect 14682 20095 15002 20096
rect 18413 19954 18479 19957
rect 22058 19954 22858 19984
rect 18413 19952 22858 19954
rect 18413 19896 18418 19952
rect 18474 19896 22858 19952
rect 18413 19894 22858 19896
rect 18413 19891 18479 19894
rect 22058 19864 22858 19894
rect 4378 19616 4698 19617
rect 4378 19552 4386 19616
rect 4450 19552 4466 19616
rect 4530 19552 4546 19616
rect 4610 19552 4626 19616
rect 4690 19552 4698 19616
rect 4378 19551 4698 19552
rect 11248 19616 11568 19617
rect 11248 19552 11256 19616
rect 11320 19552 11336 19616
rect 11400 19552 11416 19616
rect 11480 19552 11496 19616
rect 11560 19552 11568 19616
rect 11248 19551 11568 19552
rect 18117 19616 18437 19617
rect 18117 19552 18125 19616
rect 18189 19552 18205 19616
rect 18269 19552 18285 19616
rect 18349 19552 18365 19616
rect 18429 19552 18437 19616
rect 18117 19551 18437 19552
rect 7813 19072 8133 19073
rect 7813 19008 7821 19072
rect 7885 19008 7901 19072
rect 7965 19008 7981 19072
rect 8045 19008 8061 19072
rect 8125 19008 8133 19072
rect 7813 19007 8133 19008
rect 14682 19072 15002 19073
rect 14682 19008 14690 19072
rect 14754 19008 14770 19072
rect 14834 19008 14850 19072
rect 14914 19008 14930 19072
rect 14994 19008 15002 19072
rect 14682 19007 15002 19008
rect 4378 18528 4698 18529
rect 4378 18464 4386 18528
rect 4450 18464 4466 18528
rect 4530 18464 4546 18528
rect 4610 18464 4626 18528
rect 4690 18464 4698 18528
rect 4378 18463 4698 18464
rect 11248 18528 11568 18529
rect 11248 18464 11256 18528
rect 11320 18464 11336 18528
rect 11400 18464 11416 18528
rect 11480 18464 11496 18528
rect 11560 18464 11568 18528
rect 11248 18463 11568 18464
rect 18117 18528 18437 18529
rect 18117 18464 18125 18528
rect 18189 18464 18205 18528
rect 18269 18464 18285 18528
rect 18349 18464 18365 18528
rect 18429 18464 18437 18528
rect 18117 18463 18437 18464
rect 7813 17984 8133 17985
rect 7813 17920 7821 17984
rect 7885 17920 7901 17984
rect 7965 17920 7981 17984
rect 8045 17920 8061 17984
rect 8125 17920 8133 17984
rect 7813 17919 8133 17920
rect 14682 17984 15002 17985
rect 14682 17920 14690 17984
rect 14754 17920 14770 17984
rect 14834 17920 14850 17984
rect 14914 17920 14930 17984
rect 14994 17920 15002 17984
rect 14682 17919 15002 17920
rect 0 17778 800 17808
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17688 800 17718
rect 2773 17715 2839 17718
rect 4378 17440 4698 17441
rect 4378 17376 4386 17440
rect 4450 17376 4466 17440
rect 4530 17376 4546 17440
rect 4610 17376 4626 17440
rect 4690 17376 4698 17440
rect 4378 17375 4698 17376
rect 11248 17440 11568 17441
rect 11248 17376 11256 17440
rect 11320 17376 11336 17440
rect 11400 17376 11416 17440
rect 11480 17376 11496 17440
rect 11560 17376 11568 17440
rect 11248 17375 11568 17376
rect 18117 17440 18437 17441
rect 18117 17376 18125 17440
rect 18189 17376 18205 17440
rect 18269 17376 18285 17440
rect 18349 17376 18365 17440
rect 18429 17376 18437 17440
rect 18117 17375 18437 17376
rect 7813 16896 8133 16897
rect 7813 16832 7821 16896
rect 7885 16832 7901 16896
rect 7965 16832 7981 16896
rect 8045 16832 8061 16896
rect 8125 16832 8133 16896
rect 7813 16831 8133 16832
rect 14682 16896 15002 16897
rect 14682 16832 14690 16896
rect 14754 16832 14770 16896
rect 14834 16832 14850 16896
rect 14914 16832 14930 16896
rect 14994 16832 15002 16896
rect 14682 16831 15002 16832
rect 4378 16352 4698 16353
rect 4378 16288 4386 16352
rect 4450 16288 4466 16352
rect 4530 16288 4546 16352
rect 4610 16288 4626 16352
rect 4690 16288 4698 16352
rect 4378 16287 4698 16288
rect 11248 16352 11568 16353
rect 11248 16288 11256 16352
rect 11320 16288 11336 16352
rect 11400 16288 11416 16352
rect 11480 16288 11496 16352
rect 11560 16288 11568 16352
rect 11248 16287 11568 16288
rect 18117 16352 18437 16353
rect 18117 16288 18125 16352
rect 18189 16288 18205 16352
rect 18269 16288 18285 16352
rect 18349 16288 18365 16352
rect 18429 16288 18437 16352
rect 18117 16287 18437 16288
rect 7813 15808 8133 15809
rect 7813 15744 7821 15808
rect 7885 15744 7901 15808
rect 7965 15744 7981 15808
rect 8045 15744 8061 15808
rect 8125 15744 8133 15808
rect 7813 15743 8133 15744
rect 14682 15808 15002 15809
rect 14682 15744 14690 15808
rect 14754 15744 14770 15808
rect 14834 15744 14850 15808
rect 14914 15744 14930 15808
rect 14994 15744 15002 15808
rect 14682 15743 15002 15744
rect 19517 15602 19583 15605
rect 22058 15602 22858 15632
rect 19517 15600 22858 15602
rect 19517 15544 19522 15600
rect 19578 15544 22858 15600
rect 19517 15542 22858 15544
rect 19517 15539 19583 15542
rect 22058 15512 22858 15542
rect 4378 15264 4698 15265
rect 4378 15200 4386 15264
rect 4450 15200 4466 15264
rect 4530 15200 4546 15264
rect 4610 15200 4626 15264
rect 4690 15200 4698 15264
rect 4378 15199 4698 15200
rect 11248 15264 11568 15265
rect 11248 15200 11256 15264
rect 11320 15200 11336 15264
rect 11400 15200 11416 15264
rect 11480 15200 11496 15264
rect 11560 15200 11568 15264
rect 11248 15199 11568 15200
rect 18117 15264 18437 15265
rect 18117 15200 18125 15264
rect 18189 15200 18205 15264
rect 18269 15200 18285 15264
rect 18349 15200 18365 15264
rect 18429 15200 18437 15264
rect 18117 15199 18437 15200
rect 7813 14720 8133 14721
rect 7813 14656 7821 14720
rect 7885 14656 7901 14720
rect 7965 14656 7981 14720
rect 8045 14656 8061 14720
rect 8125 14656 8133 14720
rect 7813 14655 8133 14656
rect 14682 14720 15002 14721
rect 14682 14656 14690 14720
rect 14754 14656 14770 14720
rect 14834 14656 14850 14720
rect 14914 14656 14930 14720
rect 14994 14656 15002 14720
rect 14682 14655 15002 14656
rect 4378 14176 4698 14177
rect 4378 14112 4386 14176
rect 4450 14112 4466 14176
rect 4530 14112 4546 14176
rect 4610 14112 4626 14176
rect 4690 14112 4698 14176
rect 4378 14111 4698 14112
rect 11248 14176 11568 14177
rect 11248 14112 11256 14176
rect 11320 14112 11336 14176
rect 11400 14112 11416 14176
rect 11480 14112 11496 14176
rect 11560 14112 11568 14176
rect 11248 14111 11568 14112
rect 18117 14176 18437 14177
rect 18117 14112 18125 14176
rect 18189 14112 18205 14176
rect 18269 14112 18285 14176
rect 18349 14112 18365 14176
rect 18429 14112 18437 14176
rect 18117 14111 18437 14112
rect 0 13698 800 13728
rect 3417 13698 3483 13701
rect 0 13696 3483 13698
rect 0 13640 3422 13696
rect 3478 13640 3483 13696
rect 0 13638 3483 13640
rect 0 13608 800 13638
rect 3417 13635 3483 13638
rect 7813 13632 8133 13633
rect 7813 13568 7821 13632
rect 7885 13568 7901 13632
rect 7965 13568 7981 13632
rect 8045 13568 8061 13632
rect 8125 13568 8133 13632
rect 7813 13567 8133 13568
rect 14682 13632 15002 13633
rect 14682 13568 14690 13632
rect 14754 13568 14770 13632
rect 14834 13568 14850 13632
rect 14914 13568 14930 13632
rect 14994 13568 15002 13632
rect 14682 13567 15002 13568
rect 4378 13088 4698 13089
rect 4378 13024 4386 13088
rect 4450 13024 4466 13088
rect 4530 13024 4546 13088
rect 4610 13024 4626 13088
rect 4690 13024 4698 13088
rect 4378 13023 4698 13024
rect 11248 13088 11568 13089
rect 11248 13024 11256 13088
rect 11320 13024 11336 13088
rect 11400 13024 11416 13088
rect 11480 13024 11496 13088
rect 11560 13024 11568 13088
rect 11248 13023 11568 13024
rect 18117 13088 18437 13089
rect 18117 13024 18125 13088
rect 18189 13024 18205 13088
rect 18269 13024 18285 13088
rect 18349 13024 18365 13088
rect 18429 13024 18437 13088
rect 18117 13023 18437 13024
rect 7813 12544 8133 12545
rect 7813 12480 7821 12544
rect 7885 12480 7901 12544
rect 7965 12480 7981 12544
rect 8045 12480 8061 12544
rect 8125 12480 8133 12544
rect 7813 12479 8133 12480
rect 14682 12544 15002 12545
rect 14682 12480 14690 12544
rect 14754 12480 14770 12544
rect 14834 12480 14850 12544
rect 14914 12480 14930 12544
rect 14994 12480 15002 12544
rect 14682 12479 15002 12480
rect 4378 12000 4698 12001
rect 4378 11936 4386 12000
rect 4450 11936 4466 12000
rect 4530 11936 4546 12000
rect 4610 11936 4626 12000
rect 4690 11936 4698 12000
rect 4378 11935 4698 11936
rect 11248 12000 11568 12001
rect 11248 11936 11256 12000
rect 11320 11936 11336 12000
rect 11400 11936 11416 12000
rect 11480 11936 11496 12000
rect 11560 11936 11568 12000
rect 11248 11935 11568 11936
rect 18117 12000 18437 12001
rect 18117 11936 18125 12000
rect 18189 11936 18205 12000
rect 18269 11936 18285 12000
rect 18349 11936 18365 12000
rect 18429 11936 18437 12000
rect 18117 11935 18437 11936
rect 7813 11456 8133 11457
rect 7813 11392 7821 11456
rect 7885 11392 7901 11456
rect 7965 11392 7981 11456
rect 8045 11392 8061 11456
rect 8125 11392 8133 11456
rect 7813 11391 8133 11392
rect 14682 11456 15002 11457
rect 14682 11392 14690 11456
rect 14754 11392 14770 11456
rect 14834 11392 14850 11456
rect 14914 11392 14930 11456
rect 14994 11392 15002 11456
rect 14682 11391 15002 11392
rect 19701 11250 19767 11253
rect 22058 11250 22858 11280
rect 19701 11248 22858 11250
rect 19701 11192 19706 11248
rect 19762 11192 22858 11248
rect 19701 11190 22858 11192
rect 19701 11187 19767 11190
rect 22058 11160 22858 11190
rect 4378 10912 4698 10913
rect 4378 10848 4386 10912
rect 4450 10848 4466 10912
rect 4530 10848 4546 10912
rect 4610 10848 4626 10912
rect 4690 10848 4698 10912
rect 4378 10847 4698 10848
rect 11248 10912 11568 10913
rect 11248 10848 11256 10912
rect 11320 10848 11336 10912
rect 11400 10848 11416 10912
rect 11480 10848 11496 10912
rect 11560 10848 11568 10912
rect 11248 10847 11568 10848
rect 18117 10912 18437 10913
rect 18117 10848 18125 10912
rect 18189 10848 18205 10912
rect 18269 10848 18285 10912
rect 18349 10848 18365 10912
rect 18429 10848 18437 10912
rect 18117 10847 18437 10848
rect 7813 10368 8133 10369
rect 7813 10304 7821 10368
rect 7885 10304 7901 10368
rect 7965 10304 7981 10368
rect 8045 10304 8061 10368
rect 8125 10304 8133 10368
rect 7813 10303 8133 10304
rect 14682 10368 15002 10369
rect 14682 10304 14690 10368
rect 14754 10304 14770 10368
rect 14834 10304 14850 10368
rect 14914 10304 14930 10368
rect 14994 10304 15002 10368
rect 14682 10303 15002 10304
rect 4378 9824 4698 9825
rect 4378 9760 4386 9824
rect 4450 9760 4466 9824
rect 4530 9760 4546 9824
rect 4610 9760 4626 9824
rect 4690 9760 4698 9824
rect 4378 9759 4698 9760
rect 11248 9824 11568 9825
rect 11248 9760 11256 9824
rect 11320 9760 11336 9824
rect 11400 9760 11416 9824
rect 11480 9760 11496 9824
rect 11560 9760 11568 9824
rect 11248 9759 11568 9760
rect 18117 9824 18437 9825
rect 18117 9760 18125 9824
rect 18189 9760 18205 9824
rect 18269 9760 18285 9824
rect 18349 9760 18365 9824
rect 18429 9760 18437 9824
rect 18117 9759 18437 9760
rect 0 9346 800 9376
rect 4061 9346 4127 9349
rect 0 9344 4127 9346
rect 0 9288 4066 9344
rect 4122 9288 4127 9344
rect 0 9286 4127 9288
rect 0 9256 800 9286
rect 4061 9283 4127 9286
rect 7813 9280 8133 9281
rect 7813 9216 7821 9280
rect 7885 9216 7901 9280
rect 7965 9216 7981 9280
rect 8045 9216 8061 9280
rect 8125 9216 8133 9280
rect 7813 9215 8133 9216
rect 14682 9280 15002 9281
rect 14682 9216 14690 9280
rect 14754 9216 14770 9280
rect 14834 9216 14850 9280
rect 14914 9216 14930 9280
rect 14994 9216 15002 9280
rect 14682 9215 15002 9216
rect 4378 8736 4698 8737
rect 4378 8672 4386 8736
rect 4450 8672 4466 8736
rect 4530 8672 4546 8736
rect 4610 8672 4626 8736
rect 4690 8672 4698 8736
rect 4378 8671 4698 8672
rect 11248 8736 11568 8737
rect 11248 8672 11256 8736
rect 11320 8672 11336 8736
rect 11400 8672 11416 8736
rect 11480 8672 11496 8736
rect 11560 8672 11568 8736
rect 11248 8671 11568 8672
rect 18117 8736 18437 8737
rect 18117 8672 18125 8736
rect 18189 8672 18205 8736
rect 18269 8672 18285 8736
rect 18349 8672 18365 8736
rect 18429 8672 18437 8736
rect 18117 8671 18437 8672
rect 7813 8192 8133 8193
rect 7813 8128 7821 8192
rect 7885 8128 7901 8192
rect 7965 8128 7981 8192
rect 8045 8128 8061 8192
rect 8125 8128 8133 8192
rect 7813 8127 8133 8128
rect 14682 8192 15002 8193
rect 14682 8128 14690 8192
rect 14754 8128 14770 8192
rect 14834 8128 14850 8192
rect 14914 8128 14930 8192
rect 14994 8128 15002 8192
rect 14682 8127 15002 8128
rect 4378 7648 4698 7649
rect 4378 7584 4386 7648
rect 4450 7584 4466 7648
rect 4530 7584 4546 7648
rect 4610 7584 4626 7648
rect 4690 7584 4698 7648
rect 4378 7583 4698 7584
rect 11248 7648 11568 7649
rect 11248 7584 11256 7648
rect 11320 7584 11336 7648
rect 11400 7584 11416 7648
rect 11480 7584 11496 7648
rect 11560 7584 11568 7648
rect 11248 7583 11568 7584
rect 18117 7648 18437 7649
rect 18117 7584 18125 7648
rect 18189 7584 18205 7648
rect 18269 7584 18285 7648
rect 18349 7584 18365 7648
rect 18429 7584 18437 7648
rect 18117 7583 18437 7584
rect 19977 7170 20043 7173
rect 22058 7170 22858 7200
rect 19977 7168 22858 7170
rect 19977 7112 19982 7168
rect 20038 7112 22858 7168
rect 19977 7110 22858 7112
rect 19977 7107 20043 7110
rect 7813 7104 8133 7105
rect 7813 7040 7821 7104
rect 7885 7040 7901 7104
rect 7965 7040 7981 7104
rect 8045 7040 8061 7104
rect 8125 7040 8133 7104
rect 7813 7039 8133 7040
rect 14682 7104 15002 7105
rect 14682 7040 14690 7104
rect 14754 7040 14770 7104
rect 14834 7040 14850 7104
rect 14914 7040 14930 7104
rect 14994 7040 15002 7104
rect 22058 7080 22858 7110
rect 14682 7039 15002 7040
rect 4378 6560 4698 6561
rect 4378 6496 4386 6560
rect 4450 6496 4466 6560
rect 4530 6496 4546 6560
rect 4610 6496 4626 6560
rect 4690 6496 4698 6560
rect 4378 6495 4698 6496
rect 11248 6560 11568 6561
rect 11248 6496 11256 6560
rect 11320 6496 11336 6560
rect 11400 6496 11416 6560
rect 11480 6496 11496 6560
rect 11560 6496 11568 6560
rect 11248 6495 11568 6496
rect 18117 6560 18437 6561
rect 18117 6496 18125 6560
rect 18189 6496 18205 6560
rect 18269 6496 18285 6560
rect 18349 6496 18365 6560
rect 18429 6496 18437 6560
rect 18117 6495 18437 6496
rect 7813 6016 8133 6017
rect 7813 5952 7821 6016
rect 7885 5952 7901 6016
rect 7965 5952 7981 6016
rect 8045 5952 8061 6016
rect 8125 5952 8133 6016
rect 7813 5951 8133 5952
rect 14682 6016 15002 6017
rect 14682 5952 14690 6016
rect 14754 5952 14770 6016
rect 14834 5952 14850 6016
rect 14914 5952 14930 6016
rect 14994 5952 15002 6016
rect 14682 5951 15002 5952
rect 4378 5472 4698 5473
rect 4378 5408 4386 5472
rect 4450 5408 4466 5472
rect 4530 5408 4546 5472
rect 4610 5408 4626 5472
rect 4690 5408 4698 5472
rect 4378 5407 4698 5408
rect 11248 5472 11568 5473
rect 11248 5408 11256 5472
rect 11320 5408 11336 5472
rect 11400 5408 11416 5472
rect 11480 5408 11496 5472
rect 11560 5408 11568 5472
rect 11248 5407 11568 5408
rect 18117 5472 18437 5473
rect 18117 5408 18125 5472
rect 18189 5408 18205 5472
rect 18269 5408 18285 5472
rect 18349 5408 18365 5472
rect 18429 5408 18437 5472
rect 18117 5407 18437 5408
rect 0 4994 800 5024
rect 2681 4994 2747 4997
rect 0 4992 2747 4994
rect 0 4936 2686 4992
rect 2742 4936 2747 4992
rect 0 4934 2747 4936
rect 0 4904 800 4934
rect 2681 4931 2747 4934
rect 7813 4928 8133 4929
rect 7813 4864 7821 4928
rect 7885 4864 7901 4928
rect 7965 4864 7981 4928
rect 8045 4864 8061 4928
rect 8125 4864 8133 4928
rect 7813 4863 8133 4864
rect 14682 4928 15002 4929
rect 14682 4864 14690 4928
rect 14754 4864 14770 4928
rect 14834 4864 14850 4928
rect 14914 4864 14930 4928
rect 14994 4864 15002 4928
rect 14682 4863 15002 4864
rect 4378 4384 4698 4385
rect 4378 4320 4386 4384
rect 4450 4320 4466 4384
rect 4530 4320 4546 4384
rect 4610 4320 4626 4384
rect 4690 4320 4698 4384
rect 4378 4319 4698 4320
rect 11248 4384 11568 4385
rect 11248 4320 11256 4384
rect 11320 4320 11336 4384
rect 11400 4320 11416 4384
rect 11480 4320 11496 4384
rect 11560 4320 11568 4384
rect 11248 4319 11568 4320
rect 18117 4384 18437 4385
rect 18117 4320 18125 4384
rect 18189 4320 18205 4384
rect 18269 4320 18285 4384
rect 18349 4320 18365 4384
rect 18429 4320 18437 4384
rect 18117 4319 18437 4320
rect 7813 3840 8133 3841
rect 7813 3776 7821 3840
rect 7885 3776 7901 3840
rect 7965 3776 7981 3840
rect 8045 3776 8061 3840
rect 8125 3776 8133 3840
rect 7813 3775 8133 3776
rect 14682 3840 15002 3841
rect 14682 3776 14690 3840
rect 14754 3776 14770 3840
rect 14834 3776 14850 3840
rect 14914 3776 14930 3840
rect 14994 3776 15002 3840
rect 14682 3775 15002 3776
rect 4378 3296 4698 3297
rect 4378 3232 4386 3296
rect 4450 3232 4466 3296
rect 4530 3232 4546 3296
rect 4610 3232 4626 3296
rect 4690 3232 4698 3296
rect 4378 3231 4698 3232
rect 11248 3296 11568 3297
rect 11248 3232 11256 3296
rect 11320 3232 11336 3296
rect 11400 3232 11416 3296
rect 11480 3232 11496 3296
rect 11560 3232 11568 3296
rect 11248 3231 11568 3232
rect 18117 3296 18437 3297
rect 18117 3232 18125 3296
rect 18189 3232 18205 3296
rect 18269 3232 18285 3296
rect 18349 3232 18365 3296
rect 18429 3232 18437 3296
rect 18117 3231 18437 3232
rect 20345 2818 20411 2821
rect 22058 2818 22858 2848
rect 20345 2816 22858 2818
rect 20345 2760 20350 2816
rect 20406 2760 22858 2816
rect 20345 2758 22858 2760
rect 20345 2755 20411 2758
rect 7813 2752 8133 2753
rect 7813 2688 7821 2752
rect 7885 2688 7901 2752
rect 7965 2688 7981 2752
rect 8045 2688 8061 2752
rect 8125 2688 8133 2752
rect 7813 2687 8133 2688
rect 14682 2752 15002 2753
rect 14682 2688 14690 2752
rect 14754 2688 14770 2752
rect 14834 2688 14850 2752
rect 14914 2688 14930 2752
rect 14994 2688 15002 2752
rect 22058 2728 22858 2758
rect 14682 2687 15002 2688
rect 4378 2208 4698 2209
rect 4378 2144 4386 2208
rect 4450 2144 4466 2208
rect 4530 2144 4546 2208
rect 4610 2144 4626 2208
rect 4690 2144 4698 2208
rect 4378 2143 4698 2144
rect 11248 2208 11568 2209
rect 11248 2144 11256 2208
rect 11320 2144 11336 2208
rect 11400 2144 11416 2208
rect 11480 2144 11496 2208
rect 11560 2144 11568 2208
rect 11248 2143 11568 2144
rect 18117 2208 18437 2209
rect 18117 2144 18125 2208
rect 18189 2144 18205 2208
rect 18269 2144 18285 2208
rect 18349 2144 18365 2208
rect 18429 2144 18437 2208
rect 18117 2143 18437 2144
<< via3 >>
rect 7821 22332 7885 22336
rect 7821 22276 7825 22332
rect 7825 22276 7881 22332
rect 7881 22276 7885 22332
rect 7821 22272 7885 22276
rect 7901 22332 7965 22336
rect 7901 22276 7905 22332
rect 7905 22276 7961 22332
rect 7961 22276 7965 22332
rect 7901 22272 7965 22276
rect 7981 22332 8045 22336
rect 7981 22276 7985 22332
rect 7985 22276 8041 22332
rect 8041 22276 8045 22332
rect 7981 22272 8045 22276
rect 8061 22332 8125 22336
rect 8061 22276 8065 22332
rect 8065 22276 8121 22332
rect 8121 22276 8125 22332
rect 8061 22272 8125 22276
rect 14690 22332 14754 22336
rect 14690 22276 14694 22332
rect 14694 22276 14750 22332
rect 14750 22276 14754 22332
rect 14690 22272 14754 22276
rect 14770 22332 14834 22336
rect 14770 22276 14774 22332
rect 14774 22276 14830 22332
rect 14830 22276 14834 22332
rect 14770 22272 14834 22276
rect 14850 22332 14914 22336
rect 14850 22276 14854 22332
rect 14854 22276 14910 22332
rect 14910 22276 14914 22332
rect 14850 22272 14914 22276
rect 14930 22332 14994 22336
rect 14930 22276 14934 22332
rect 14934 22276 14990 22332
rect 14990 22276 14994 22332
rect 14930 22272 14994 22276
rect 4386 21788 4450 21792
rect 4386 21732 4390 21788
rect 4390 21732 4446 21788
rect 4446 21732 4450 21788
rect 4386 21728 4450 21732
rect 4466 21788 4530 21792
rect 4466 21732 4470 21788
rect 4470 21732 4526 21788
rect 4526 21732 4530 21788
rect 4466 21728 4530 21732
rect 4546 21788 4610 21792
rect 4546 21732 4550 21788
rect 4550 21732 4606 21788
rect 4606 21732 4610 21788
rect 4546 21728 4610 21732
rect 4626 21788 4690 21792
rect 4626 21732 4630 21788
rect 4630 21732 4686 21788
rect 4686 21732 4690 21788
rect 4626 21728 4690 21732
rect 11256 21788 11320 21792
rect 11256 21732 11260 21788
rect 11260 21732 11316 21788
rect 11316 21732 11320 21788
rect 11256 21728 11320 21732
rect 11336 21788 11400 21792
rect 11336 21732 11340 21788
rect 11340 21732 11396 21788
rect 11396 21732 11400 21788
rect 11336 21728 11400 21732
rect 11416 21788 11480 21792
rect 11416 21732 11420 21788
rect 11420 21732 11476 21788
rect 11476 21732 11480 21788
rect 11416 21728 11480 21732
rect 11496 21788 11560 21792
rect 11496 21732 11500 21788
rect 11500 21732 11556 21788
rect 11556 21732 11560 21788
rect 11496 21728 11560 21732
rect 18125 21788 18189 21792
rect 18125 21732 18129 21788
rect 18129 21732 18185 21788
rect 18185 21732 18189 21788
rect 18125 21728 18189 21732
rect 18205 21788 18269 21792
rect 18205 21732 18209 21788
rect 18209 21732 18265 21788
rect 18265 21732 18269 21788
rect 18205 21728 18269 21732
rect 18285 21788 18349 21792
rect 18285 21732 18289 21788
rect 18289 21732 18345 21788
rect 18345 21732 18349 21788
rect 18285 21728 18349 21732
rect 18365 21788 18429 21792
rect 18365 21732 18369 21788
rect 18369 21732 18425 21788
rect 18425 21732 18429 21788
rect 18365 21728 18429 21732
rect 7821 21244 7885 21248
rect 7821 21188 7825 21244
rect 7825 21188 7881 21244
rect 7881 21188 7885 21244
rect 7821 21184 7885 21188
rect 7901 21244 7965 21248
rect 7901 21188 7905 21244
rect 7905 21188 7961 21244
rect 7961 21188 7965 21244
rect 7901 21184 7965 21188
rect 7981 21244 8045 21248
rect 7981 21188 7985 21244
rect 7985 21188 8041 21244
rect 8041 21188 8045 21244
rect 7981 21184 8045 21188
rect 8061 21244 8125 21248
rect 8061 21188 8065 21244
rect 8065 21188 8121 21244
rect 8121 21188 8125 21244
rect 8061 21184 8125 21188
rect 14690 21244 14754 21248
rect 14690 21188 14694 21244
rect 14694 21188 14750 21244
rect 14750 21188 14754 21244
rect 14690 21184 14754 21188
rect 14770 21244 14834 21248
rect 14770 21188 14774 21244
rect 14774 21188 14830 21244
rect 14830 21188 14834 21244
rect 14770 21184 14834 21188
rect 14850 21244 14914 21248
rect 14850 21188 14854 21244
rect 14854 21188 14910 21244
rect 14910 21188 14914 21244
rect 14850 21184 14914 21188
rect 14930 21244 14994 21248
rect 14930 21188 14934 21244
rect 14934 21188 14990 21244
rect 14990 21188 14994 21244
rect 14930 21184 14994 21188
rect 4386 20700 4450 20704
rect 4386 20644 4390 20700
rect 4390 20644 4446 20700
rect 4446 20644 4450 20700
rect 4386 20640 4450 20644
rect 4466 20700 4530 20704
rect 4466 20644 4470 20700
rect 4470 20644 4526 20700
rect 4526 20644 4530 20700
rect 4466 20640 4530 20644
rect 4546 20700 4610 20704
rect 4546 20644 4550 20700
rect 4550 20644 4606 20700
rect 4606 20644 4610 20700
rect 4546 20640 4610 20644
rect 4626 20700 4690 20704
rect 4626 20644 4630 20700
rect 4630 20644 4686 20700
rect 4686 20644 4690 20700
rect 4626 20640 4690 20644
rect 11256 20700 11320 20704
rect 11256 20644 11260 20700
rect 11260 20644 11316 20700
rect 11316 20644 11320 20700
rect 11256 20640 11320 20644
rect 11336 20700 11400 20704
rect 11336 20644 11340 20700
rect 11340 20644 11396 20700
rect 11396 20644 11400 20700
rect 11336 20640 11400 20644
rect 11416 20700 11480 20704
rect 11416 20644 11420 20700
rect 11420 20644 11476 20700
rect 11476 20644 11480 20700
rect 11416 20640 11480 20644
rect 11496 20700 11560 20704
rect 11496 20644 11500 20700
rect 11500 20644 11556 20700
rect 11556 20644 11560 20700
rect 11496 20640 11560 20644
rect 18125 20700 18189 20704
rect 18125 20644 18129 20700
rect 18129 20644 18185 20700
rect 18185 20644 18189 20700
rect 18125 20640 18189 20644
rect 18205 20700 18269 20704
rect 18205 20644 18209 20700
rect 18209 20644 18265 20700
rect 18265 20644 18269 20700
rect 18205 20640 18269 20644
rect 18285 20700 18349 20704
rect 18285 20644 18289 20700
rect 18289 20644 18345 20700
rect 18345 20644 18349 20700
rect 18285 20640 18349 20644
rect 18365 20700 18429 20704
rect 18365 20644 18369 20700
rect 18369 20644 18425 20700
rect 18425 20644 18429 20700
rect 18365 20640 18429 20644
rect 7821 20156 7885 20160
rect 7821 20100 7825 20156
rect 7825 20100 7881 20156
rect 7881 20100 7885 20156
rect 7821 20096 7885 20100
rect 7901 20156 7965 20160
rect 7901 20100 7905 20156
rect 7905 20100 7961 20156
rect 7961 20100 7965 20156
rect 7901 20096 7965 20100
rect 7981 20156 8045 20160
rect 7981 20100 7985 20156
rect 7985 20100 8041 20156
rect 8041 20100 8045 20156
rect 7981 20096 8045 20100
rect 8061 20156 8125 20160
rect 8061 20100 8065 20156
rect 8065 20100 8121 20156
rect 8121 20100 8125 20156
rect 8061 20096 8125 20100
rect 14690 20156 14754 20160
rect 14690 20100 14694 20156
rect 14694 20100 14750 20156
rect 14750 20100 14754 20156
rect 14690 20096 14754 20100
rect 14770 20156 14834 20160
rect 14770 20100 14774 20156
rect 14774 20100 14830 20156
rect 14830 20100 14834 20156
rect 14770 20096 14834 20100
rect 14850 20156 14914 20160
rect 14850 20100 14854 20156
rect 14854 20100 14910 20156
rect 14910 20100 14914 20156
rect 14850 20096 14914 20100
rect 14930 20156 14994 20160
rect 14930 20100 14934 20156
rect 14934 20100 14990 20156
rect 14990 20100 14994 20156
rect 14930 20096 14994 20100
rect 4386 19612 4450 19616
rect 4386 19556 4390 19612
rect 4390 19556 4446 19612
rect 4446 19556 4450 19612
rect 4386 19552 4450 19556
rect 4466 19612 4530 19616
rect 4466 19556 4470 19612
rect 4470 19556 4526 19612
rect 4526 19556 4530 19612
rect 4466 19552 4530 19556
rect 4546 19612 4610 19616
rect 4546 19556 4550 19612
rect 4550 19556 4606 19612
rect 4606 19556 4610 19612
rect 4546 19552 4610 19556
rect 4626 19612 4690 19616
rect 4626 19556 4630 19612
rect 4630 19556 4686 19612
rect 4686 19556 4690 19612
rect 4626 19552 4690 19556
rect 11256 19612 11320 19616
rect 11256 19556 11260 19612
rect 11260 19556 11316 19612
rect 11316 19556 11320 19612
rect 11256 19552 11320 19556
rect 11336 19612 11400 19616
rect 11336 19556 11340 19612
rect 11340 19556 11396 19612
rect 11396 19556 11400 19612
rect 11336 19552 11400 19556
rect 11416 19612 11480 19616
rect 11416 19556 11420 19612
rect 11420 19556 11476 19612
rect 11476 19556 11480 19612
rect 11416 19552 11480 19556
rect 11496 19612 11560 19616
rect 11496 19556 11500 19612
rect 11500 19556 11556 19612
rect 11556 19556 11560 19612
rect 11496 19552 11560 19556
rect 18125 19612 18189 19616
rect 18125 19556 18129 19612
rect 18129 19556 18185 19612
rect 18185 19556 18189 19612
rect 18125 19552 18189 19556
rect 18205 19612 18269 19616
rect 18205 19556 18209 19612
rect 18209 19556 18265 19612
rect 18265 19556 18269 19612
rect 18205 19552 18269 19556
rect 18285 19612 18349 19616
rect 18285 19556 18289 19612
rect 18289 19556 18345 19612
rect 18345 19556 18349 19612
rect 18285 19552 18349 19556
rect 18365 19612 18429 19616
rect 18365 19556 18369 19612
rect 18369 19556 18425 19612
rect 18425 19556 18429 19612
rect 18365 19552 18429 19556
rect 7821 19068 7885 19072
rect 7821 19012 7825 19068
rect 7825 19012 7881 19068
rect 7881 19012 7885 19068
rect 7821 19008 7885 19012
rect 7901 19068 7965 19072
rect 7901 19012 7905 19068
rect 7905 19012 7961 19068
rect 7961 19012 7965 19068
rect 7901 19008 7965 19012
rect 7981 19068 8045 19072
rect 7981 19012 7985 19068
rect 7985 19012 8041 19068
rect 8041 19012 8045 19068
rect 7981 19008 8045 19012
rect 8061 19068 8125 19072
rect 8061 19012 8065 19068
rect 8065 19012 8121 19068
rect 8121 19012 8125 19068
rect 8061 19008 8125 19012
rect 14690 19068 14754 19072
rect 14690 19012 14694 19068
rect 14694 19012 14750 19068
rect 14750 19012 14754 19068
rect 14690 19008 14754 19012
rect 14770 19068 14834 19072
rect 14770 19012 14774 19068
rect 14774 19012 14830 19068
rect 14830 19012 14834 19068
rect 14770 19008 14834 19012
rect 14850 19068 14914 19072
rect 14850 19012 14854 19068
rect 14854 19012 14910 19068
rect 14910 19012 14914 19068
rect 14850 19008 14914 19012
rect 14930 19068 14994 19072
rect 14930 19012 14934 19068
rect 14934 19012 14990 19068
rect 14990 19012 14994 19068
rect 14930 19008 14994 19012
rect 4386 18524 4450 18528
rect 4386 18468 4390 18524
rect 4390 18468 4446 18524
rect 4446 18468 4450 18524
rect 4386 18464 4450 18468
rect 4466 18524 4530 18528
rect 4466 18468 4470 18524
rect 4470 18468 4526 18524
rect 4526 18468 4530 18524
rect 4466 18464 4530 18468
rect 4546 18524 4610 18528
rect 4546 18468 4550 18524
rect 4550 18468 4606 18524
rect 4606 18468 4610 18524
rect 4546 18464 4610 18468
rect 4626 18524 4690 18528
rect 4626 18468 4630 18524
rect 4630 18468 4686 18524
rect 4686 18468 4690 18524
rect 4626 18464 4690 18468
rect 11256 18524 11320 18528
rect 11256 18468 11260 18524
rect 11260 18468 11316 18524
rect 11316 18468 11320 18524
rect 11256 18464 11320 18468
rect 11336 18524 11400 18528
rect 11336 18468 11340 18524
rect 11340 18468 11396 18524
rect 11396 18468 11400 18524
rect 11336 18464 11400 18468
rect 11416 18524 11480 18528
rect 11416 18468 11420 18524
rect 11420 18468 11476 18524
rect 11476 18468 11480 18524
rect 11416 18464 11480 18468
rect 11496 18524 11560 18528
rect 11496 18468 11500 18524
rect 11500 18468 11556 18524
rect 11556 18468 11560 18524
rect 11496 18464 11560 18468
rect 18125 18524 18189 18528
rect 18125 18468 18129 18524
rect 18129 18468 18185 18524
rect 18185 18468 18189 18524
rect 18125 18464 18189 18468
rect 18205 18524 18269 18528
rect 18205 18468 18209 18524
rect 18209 18468 18265 18524
rect 18265 18468 18269 18524
rect 18205 18464 18269 18468
rect 18285 18524 18349 18528
rect 18285 18468 18289 18524
rect 18289 18468 18345 18524
rect 18345 18468 18349 18524
rect 18285 18464 18349 18468
rect 18365 18524 18429 18528
rect 18365 18468 18369 18524
rect 18369 18468 18425 18524
rect 18425 18468 18429 18524
rect 18365 18464 18429 18468
rect 7821 17980 7885 17984
rect 7821 17924 7825 17980
rect 7825 17924 7881 17980
rect 7881 17924 7885 17980
rect 7821 17920 7885 17924
rect 7901 17980 7965 17984
rect 7901 17924 7905 17980
rect 7905 17924 7961 17980
rect 7961 17924 7965 17980
rect 7901 17920 7965 17924
rect 7981 17980 8045 17984
rect 7981 17924 7985 17980
rect 7985 17924 8041 17980
rect 8041 17924 8045 17980
rect 7981 17920 8045 17924
rect 8061 17980 8125 17984
rect 8061 17924 8065 17980
rect 8065 17924 8121 17980
rect 8121 17924 8125 17980
rect 8061 17920 8125 17924
rect 14690 17980 14754 17984
rect 14690 17924 14694 17980
rect 14694 17924 14750 17980
rect 14750 17924 14754 17980
rect 14690 17920 14754 17924
rect 14770 17980 14834 17984
rect 14770 17924 14774 17980
rect 14774 17924 14830 17980
rect 14830 17924 14834 17980
rect 14770 17920 14834 17924
rect 14850 17980 14914 17984
rect 14850 17924 14854 17980
rect 14854 17924 14910 17980
rect 14910 17924 14914 17980
rect 14850 17920 14914 17924
rect 14930 17980 14994 17984
rect 14930 17924 14934 17980
rect 14934 17924 14990 17980
rect 14990 17924 14994 17980
rect 14930 17920 14994 17924
rect 4386 17436 4450 17440
rect 4386 17380 4390 17436
rect 4390 17380 4446 17436
rect 4446 17380 4450 17436
rect 4386 17376 4450 17380
rect 4466 17436 4530 17440
rect 4466 17380 4470 17436
rect 4470 17380 4526 17436
rect 4526 17380 4530 17436
rect 4466 17376 4530 17380
rect 4546 17436 4610 17440
rect 4546 17380 4550 17436
rect 4550 17380 4606 17436
rect 4606 17380 4610 17436
rect 4546 17376 4610 17380
rect 4626 17436 4690 17440
rect 4626 17380 4630 17436
rect 4630 17380 4686 17436
rect 4686 17380 4690 17436
rect 4626 17376 4690 17380
rect 11256 17436 11320 17440
rect 11256 17380 11260 17436
rect 11260 17380 11316 17436
rect 11316 17380 11320 17436
rect 11256 17376 11320 17380
rect 11336 17436 11400 17440
rect 11336 17380 11340 17436
rect 11340 17380 11396 17436
rect 11396 17380 11400 17436
rect 11336 17376 11400 17380
rect 11416 17436 11480 17440
rect 11416 17380 11420 17436
rect 11420 17380 11476 17436
rect 11476 17380 11480 17436
rect 11416 17376 11480 17380
rect 11496 17436 11560 17440
rect 11496 17380 11500 17436
rect 11500 17380 11556 17436
rect 11556 17380 11560 17436
rect 11496 17376 11560 17380
rect 18125 17436 18189 17440
rect 18125 17380 18129 17436
rect 18129 17380 18185 17436
rect 18185 17380 18189 17436
rect 18125 17376 18189 17380
rect 18205 17436 18269 17440
rect 18205 17380 18209 17436
rect 18209 17380 18265 17436
rect 18265 17380 18269 17436
rect 18205 17376 18269 17380
rect 18285 17436 18349 17440
rect 18285 17380 18289 17436
rect 18289 17380 18345 17436
rect 18345 17380 18349 17436
rect 18285 17376 18349 17380
rect 18365 17436 18429 17440
rect 18365 17380 18369 17436
rect 18369 17380 18425 17436
rect 18425 17380 18429 17436
rect 18365 17376 18429 17380
rect 7821 16892 7885 16896
rect 7821 16836 7825 16892
rect 7825 16836 7881 16892
rect 7881 16836 7885 16892
rect 7821 16832 7885 16836
rect 7901 16892 7965 16896
rect 7901 16836 7905 16892
rect 7905 16836 7961 16892
rect 7961 16836 7965 16892
rect 7901 16832 7965 16836
rect 7981 16892 8045 16896
rect 7981 16836 7985 16892
rect 7985 16836 8041 16892
rect 8041 16836 8045 16892
rect 7981 16832 8045 16836
rect 8061 16892 8125 16896
rect 8061 16836 8065 16892
rect 8065 16836 8121 16892
rect 8121 16836 8125 16892
rect 8061 16832 8125 16836
rect 14690 16892 14754 16896
rect 14690 16836 14694 16892
rect 14694 16836 14750 16892
rect 14750 16836 14754 16892
rect 14690 16832 14754 16836
rect 14770 16892 14834 16896
rect 14770 16836 14774 16892
rect 14774 16836 14830 16892
rect 14830 16836 14834 16892
rect 14770 16832 14834 16836
rect 14850 16892 14914 16896
rect 14850 16836 14854 16892
rect 14854 16836 14910 16892
rect 14910 16836 14914 16892
rect 14850 16832 14914 16836
rect 14930 16892 14994 16896
rect 14930 16836 14934 16892
rect 14934 16836 14990 16892
rect 14990 16836 14994 16892
rect 14930 16832 14994 16836
rect 4386 16348 4450 16352
rect 4386 16292 4390 16348
rect 4390 16292 4446 16348
rect 4446 16292 4450 16348
rect 4386 16288 4450 16292
rect 4466 16348 4530 16352
rect 4466 16292 4470 16348
rect 4470 16292 4526 16348
rect 4526 16292 4530 16348
rect 4466 16288 4530 16292
rect 4546 16348 4610 16352
rect 4546 16292 4550 16348
rect 4550 16292 4606 16348
rect 4606 16292 4610 16348
rect 4546 16288 4610 16292
rect 4626 16348 4690 16352
rect 4626 16292 4630 16348
rect 4630 16292 4686 16348
rect 4686 16292 4690 16348
rect 4626 16288 4690 16292
rect 11256 16348 11320 16352
rect 11256 16292 11260 16348
rect 11260 16292 11316 16348
rect 11316 16292 11320 16348
rect 11256 16288 11320 16292
rect 11336 16348 11400 16352
rect 11336 16292 11340 16348
rect 11340 16292 11396 16348
rect 11396 16292 11400 16348
rect 11336 16288 11400 16292
rect 11416 16348 11480 16352
rect 11416 16292 11420 16348
rect 11420 16292 11476 16348
rect 11476 16292 11480 16348
rect 11416 16288 11480 16292
rect 11496 16348 11560 16352
rect 11496 16292 11500 16348
rect 11500 16292 11556 16348
rect 11556 16292 11560 16348
rect 11496 16288 11560 16292
rect 18125 16348 18189 16352
rect 18125 16292 18129 16348
rect 18129 16292 18185 16348
rect 18185 16292 18189 16348
rect 18125 16288 18189 16292
rect 18205 16348 18269 16352
rect 18205 16292 18209 16348
rect 18209 16292 18265 16348
rect 18265 16292 18269 16348
rect 18205 16288 18269 16292
rect 18285 16348 18349 16352
rect 18285 16292 18289 16348
rect 18289 16292 18345 16348
rect 18345 16292 18349 16348
rect 18285 16288 18349 16292
rect 18365 16348 18429 16352
rect 18365 16292 18369 16348
rect 18369 16292 18425 16348
rect 18425 16292 18429 16348
rect 18365 16288 18429 16292
rect 7821 15804 7885 15808
rect 7821 15748 7825 15804
rect 7825 15748 7881 15804
rect 7881 15748 7885 15804
rect 7821 15744 7885 15748
rect 7901 15804 7965 15808
rect 7901 15748 7905 15804
rect 7905 15748 7961 15804
rect 7961 15748 7965 15804
rect 7901 15744 7965 15748
rect 7981 15804 8045 15808
rect 7981 15748 7985 15804
rect 7985 15748 8041 15804
rect 8041 15748 8045 15804
rect 7981 15744 8045 15748
rect 8061 15804 8125 15808
rect 8061 15748 8065 15804
rect 8065 15748 8121 15804
rect 8121 15748 8125 15804
rect 8061 15744 8125 15748
rect 14690 15804 14754 15808
rect 14690 15748 14694 15804
rect 14694 15748 14750 15804
rect 14750 15748 14754 15804
rect 14690 15744 14754 15748
rect 14770 15804 14834 15808
rect 14770 15748 14774 15804
rect 14774 15748 14830 15804
rect 14830 15748 14834 15804
rect 14770 15744 14834 15748
rect 14850 15804 14914 15808
rect 14850 15748 14854 15804
rect 14854 15748 14910 15804
rect 14910 15748 14914 15804
rect 14850 15744 14914 15748
rect 14930 15804 14994 15808
rect 14930 15748 14934 15804
rect 14934 15748 14990 15804
rect 14990 15748 14994 15804
rect 14930 15744 14994 15748
rect 4386 15260 4450 15264
rect 4386 15204 4390 15260
rect 4390 15204 4446 15260
rect 4446 15204 4450 15260
rect 4386 15200 4450 15204
rect 4466 15260 4530 15264
rect 4466 15204 4470 15260
rect 4470 15204 4526 15260
rect 4526 15204 4530 15260
rect 4466 15200 4530 15204
rect 4546 15260 4610 15264
rect 4546 15204 4550 15260
rect 4550 15204 4606 15260
rect 4606 15204 4610 15260
rect 4546 15200 4610 15204
rect 4626 15260 4690 15264
rect 4626 15204 4630 15260
rect 4630 15204 4686 15260
rect 4686 15204 4690 15260
rect 4626 15200 4690 15204
rect 11256 15260 11320 15264
rect 11256 15204 11260 15260
rect 11260 15204 11316 15260
rect 11316 15204 11320 15260
rect 11256 15200 11320 15204
rect 11336 15260 11400 15264
rect 11336 15204 11340 15260
rect 11340 15204 11396 15260
rect 11396 15204 11400 15260
rect 11336 15200 11400 15204
rect 11416 15260 11480 15264
rect 11416 15204 11420 15260
rect 11420 15204 11476 15260
rect 11476 15204 11480 15260
rect 11416 15200 11480 15204
rect 11496 15260 11560 15264
rect 11496 15204 11500 15260
rect 11500 15204 11556 15260
rect 11556 15204 11560 15260
rect 11496 15200 11560 15204
rect 18125 15260 18189 15264
rect 18125 15204 18129 15260
rect 18129 15204 18185 15260
rect 18185 15204 18189 15260
rect 18125 15200 18189 15204
rect 18205 15260 18269 15264
rect 18205 15204 18209 15260
rect 18209 15204 18265 15260
rect 18265 15204 18269 15260
rect 18205 15200 18269 15204
rect 18285 15260 18349 15264
rect 18285 15204 18289 15260
rect 18289 15204 18345 15260
rect 18345 15204 18349 15260
rect 18285 15200 18349 15204
rect 18365 15260 18429 15264
rect 18365 15204 18369 15260
rect 18369 15204 18425 15260
rect 18425 15204 18429 15260
rect 18365 15200 18429 15204
rect 7821 14716 7885 14720
rect 7821 14660 7825 14716
rect 7825 14660 7881 14716
rect 7881 14660 7885 14716
rect 7821 14656 7885 14660
rect 7901 14716 7965 14720
rect 7901 14660 7905 14716
rect 7905 14660 7961 14716
rect 7961 14660 7965 14716
rect 7901 14656 7965 14660
rect 7981 14716 8045 14720
rect 7981 14660 7985 14716
rect 7985 14660 8041 14716
rect 8041 14660 8045 14716
rect 7981 14656 8045 14660
rect 8061 14716 8125 14720
rect 8061 14660 8065 14716
rect 8065 14660 8121 14716
rect 8121 14660 8125 14716
rect 8061 14656 8125 14660
rect 14690 14716 14754 14720
rect 14690 14660 14694 14716
rect 14694 14660 14750 14716
rect 14750 14660 14754 14716
rect 14690 14656 14754 14660
rect 14770 14716 14834 14720
rect 14770 14660 14774 14716
rect 14774 14660 14830 14716
rect 14830 14660 14834 14716
rect 14770 14656 14834 14660
rect 14850 14716 14914 14720
rect 14850 14660 14854 14716
rect 14854 14660 14910 14716
rect 14910 14660 14914 14716
rect 14850 14656 14914 14660
rect 14930 14716 14994 14720
rect 14930 14660 14934 14716
rect 14934 14660 14990 14716
rect 14990 14660 14994 14716
rect 14930 14656 14994 14660
rect 4386 14172 4450 14176
rect 4386 14116 4390 14172
rect 4390 14116 4446 14172
rect 4446 14116 4450 14172
rect 4386 14112 4450 14116
rect 4466 14172 4530 14176
rect 4466 14116 4470 14172
rect 4470 14116 4526 14172
rect 4526 14116 4530 14172
rect 4466 14112 4530 14116
rect 4546 14172 4610 14176
rect 4546 14116 4550 14172
rect 4550 14116 4606 14172
rect 4606 14116 4610 14172
rect 4546 14112 4610 14116
rect 4626 14172 4690 14176
rect 4626 14116 4630 14172
rect 4630 14116 4686 14172
rect 4686 14116 4690 14172
rect 4626 14112 4690 14116
rect 11256 14172 11320 14176
rect 11256 14116 11260 14172
rect 11260 14116 11316 14172
rect 11316 14116 11320 14172
rect 11256 14112 11320 14116
rect 11336 14172 11400 14176
rect 11336 14116 11340 14172
rect 11340 14116 11396 14172
rect 11396 14116 11400 14172
rect 11336 14112 11400 14116
rect 11416 14172 11480 14176
rect 11416 14116 11420 14172
rect 11420 14116 11476 14172
rect 11476 14116 11480 14172
rect 11416 14112 11480 14116
rect 11496 14172 11560 14176
rect 11496 14116 11500 14172
rect 11500 14116 11556 14172
rect 11556 14116 11560 14172
rect 11496 14112 11560 14116
rect 18125 14172 18189 14176
rect 18125 14116 18129 14172
rect 18129 14116 18185 14172
rect 18185 14116 18189 14172
rect 18125 14112 18189 14116
rect 18205 14172 18269 14176
rect 18205 14116 18209 14172
rect 18209 14116 18265 14172
rect 18265 14116 18269 14172
rect 18205 14112 18269 14116
rect 18285 14172 18349 14176
rect 18285 14116 18289 14172
rect 18289 14116 18345 14172
rect 18345 14116 18349 14172
rect 18285 14112 18349 14116
rect 18365 14172 18429 14176
rect 18365 14116 18369 14172
rect 18369 14116 18425 14172
rect 18425 14116 18429 14172
rect 18365 14112 18429 14116
rect 7821 13628 7885 13632
rect 7821 13572 7825 13628
rect 7825 13572 7881 13628
rect 7881 13572 7885 13628
rect 7821 13568 7885 13572
rect 7901 13628 7965 13632
rect 7901 13572 7905 13628
rect 7905 13572 7961 13628
rect 7961 13572 7965 13628
rect 7901 13568 7965 13572
rect 7981 13628 8045 13632
rect 7981 13572 7985 13628
rect 7985 13572 8041 13628
rect 8041 13572 8045 13628
rect 7981 13568 8045 13572
rect 8061 13628 8125 13632
rect 8061 13572 8065 13628
rect 8065 13572 8121 13628
rect 8121 13572 8125 13628
rect 8061 13568 8125 13572
rect 14690 13628 14754 13632
rect 14690 13572 14694 13628
rect 14694 13572 14750 13628
rect 14750 13572 14754 13628
rect 14690 13568 14754 13572
rect 14770 13628 14834 13632
rect 14770 13572 14774 13628
rect 14774 13572 14830 13628
rect 14830 13572 14834 13628
rect 14770 13568 14834 13572
rect 14850 13628 14914 13632
rect 14850 13572 14854 13628
rect 14854 13572 14910 13628
rect 14910 13572 14914 13628
rect 14850 13568 14914 13572
rect 14930 13628 14994 13632
rect 14930 13572 14934 13628
rect 14934 13572 14990 13628
rect 14990 13572 14994 13628
rect 14930 13568 14994 13572
rect 4386 13084 4450 13088
rect 4386 13028 4390 13084
rect 4390 13028 4446 13084
rect 4446 13028 4450 13084
rect 4386 13024 4450 13028
rect 4466 13084 4530 13088
rect 4466 13028 4470 13084
rect 4470 13028 4526 13084
rect 4526 13028 4530 13084
rect 4466 13024 4530 13028
rect 4546 13084 4610 13088
rect 4546 13028 4550 13084
rect 4550 13028 4606 13084
rect 4606 13028 4610 13084
rect 4546 13024 4610 13028
rect 4626 13084 4690 13088
rect 4626 13028 4630 13084
rect 4630 13028 4686 13084
rect 4686 13028 4690 13084
rect 4626 13024 4690 13028
rect 11256 13084 11320 13088
rect 11256 13028 11260 13084
rect 11260 13028 11316 13084
rect 11316 13028 11320 13084
rect 11256 13024 11320 13028
rect 11336 13084 11400 13088
rect 11336 13028 11340 13084
rect 11340 13028 11396 13084
rect 11396 13028 11400 13084
rect 11336 13024 11400 13028
rect 11416 13084 11480 13088
rect 11416 13028 11420 13084
rect 11420 13028 11476 13084
rect 11476 13028 11480 13084
rect 11416 13024 11480 13028
rect 11496 13084 11560 13088
rect 11496 13028 11500 13084
rect 11500 13028 11556 13084
rect 11556 13028 11560 13084
rect 11496 13024 11560 13028
rect 18125 13084 18189 13088
rect 18125 13028 18129 13084
rect 18129 13028 18185 13084
rect 18185 13028 18189 13084
rect 18125 13024 18189 13028
rect 18205 13084 18269 13088
rect 18205 13028 18209 13084
rect 18209 13028 18265 13084
rect 18265 13028 18269 13084
rect 18205 13024 18269 13028
rect 18285 13084 18349 13088
rect 18285 13028 18289 13084
rect 18289 13028 18345 13084
rect 18345 13028 18349 13084
rect 18285 13024 18349 13028
rect 18365 13084 18429 13088
rect 18365 13028 18369 13084
rect 18369 13028 18425 13084
rect 18425 13028 18429 13084
rect 18365 13024 18429 13028
rect 7821 12540 7885 12544
rect 7821 12484 7825 12540
rect 7825 12484 7881 12540
rect 7881 12484 7885 12540
rect 7821 12480 7885 12484
rect 7901 12540 7965 12544
rect 7901 12484 7905 12540
rect 7905 12484 7961 12540
rect 7961 12484 7965 12540
rect 7901 12480 7965 12484
rect 7981 12540 8045 12544
rect 7981 12484 7985 12540
rect 7985 12484 8041 12540
rect 8041 12484 8045 12540
rect 7981 12480 8045 12484
rect 8061 12540 8125 12544
rect 8061 12484 8065 12540
rect 8065 12484 8121 12540
rect 8121 12484 8125 12540
rect 8061 12480 8125 12484
rect 14690 12540 14754 12544
rect 14690 12484 14694 12540
rect 14694 12484 14750 12540
rect 14750 12484 14754 12540
rect 14690 12480 14754 12484
rect 14770 12540 14834 12544
rect 14770 12484 14774 12540
rect 14774 12484 14830 12540
rect 14830 12484 14834 12540
rect 14770 12480 14834 12484
rect 14850 12540 14914 12544
rect 14850 12484 14854 12540
rect 14854 12484 14910 12540
rect 14910 12484 14914 12540
rect 14850 12480 14914 12484
rect 14930 12540 14994 12544
rect 14930 12484 14934 12540
rect 14934 12484 14990 12540
rect 14990 12484 14994 12540
rect 14930 12480 14994 12484
rect 4386 11996 4450 12000
rect 4386 11940 4390 11996
rect 4390 11940 4446 11996
rect 4446 11940 4450 11996
rect 4386 11936 4450 11940
rect 4466 11996 4530 12000
rect 4466 11940 4470 11996
rect 4470 11940 4526 11996
rect 4526 11940 4530 11996
rect 4466 11936 4530 11940
rect 4546 11996 4610 12000
rect 4546 11940 4550 11996
rect 4550 11940 4606 11996
rect 4606 11940 4610 11996
rect 4546 11936 4610 11940
rect 4626 11996 4690 12000
rect 4626 11940 4630 11996
rect 4630 11940 4686 11996
rect 4686 11940 4690 11996
rect 4626 11936 4690 11940
rect 11256 11996 11320 12000
rect 11256 11940 11260 11996
rect 11260 11940 11316 11996
rect 11316 11940 11320 11996
rect 11256 11936 11320 11940
rect 11336 11996 11400 12000
rect 11336 11940 11340 11996
rect 11340 11940 11396 11996
rect 11396 11940 11400 11996
rect 11336 11936 11400 11940
rect 11416 11996 11480 12000
rect 11416 11940 11420 11996
rect 11420 11940 11476 11996
rect 11476 11940 11480 11996
rect 11416 11936 11480 11940
rect 11496 11996 11560 12000
rect 11496 11940 11500 11996
rect 11500 11940 11556 11996
rect 11556 11940 11560 11996
rect 11496 11936 11560 11940
rect 18125 11996 18189 12000
rect 18125 11940 18129 11996
rect 18129 11940 18185 11996
rect 18185 11940 18189 11996
rect 18125 11936 18189 11940
rect 18205 11996 18269 12000
rect 18205 11940 18209 11996
rect 18209 11940 18265 11996
rect 18265 11940 18269 11996
rect 18205 11936 18269 11940
rect 18285 11996 18349 12000
rect 18285 11940 18289 11996
rect 18289 11940 18345 11996
rect 18345 11940 18349 11996
rect 18285 11936 18349 11940
rect 18365 11996 18429 12000
rect 18365 11940 18369 11996
rect 18369 11940 18425 11996
rect 18425 11940 18429 11996
rect 18365 11936 18429 11940
rect 7821 11452 7885 11456
rect 7821 11396 7825 11452
rect 7825 11396 7881 11452
rect 7881 11396 7885 11452
rect 7821 11392 7885 11396
rect 7901 11452 7965 11456
rect 7901 11396 7905 11452
rect 7905 11396 7961 11452
rect 7961 11396 7965 11452
rect 7901 11392 7965 11396
rect 7981 11452 8045 11456
rect 7981 11396 7985 11452
rect 7985 11396 8041 11452
rect 8041 11396 8045 11452
rect 7981 11392 8045 11396
rect 8061 11452 8125 11456
rect 8061 11396 8065 11452
rect 8065 11396 8121 11452
rect 8121 11396 8125 11452
rect 8061 11392 8125 11396
rect 14690 11452 14754 11456
rect 14690 11396 14694 11452
rect 14694 11396 14750 11452
rect 14750 11396 14754 11452
rect 14690 11392 14754 11396
rect 14770 11452 14834 11456
rect 14770 11396 14774 11452
rect 14774 11396 14830 11452
rect 14830 11396 14834 11452
rect 14770 11392 14834 11396
rect 14850 11452 14914 11456
rect 14850 11396 14854 11452
rect 14854 11396 14910 11452
rect 14910 11396 14914 11452
rect 14850 11392 14914 11396
rect 14930 11452 14994 11456
rect 14930 11396 14934 11452
rect 14934 11396 14990 11452
rect 14990 11396 14994 11452
rect 14930 11392 14994 11396
rect 4386 10908 4450 10912
rect 4386 10852 4390 10908
rect 4390 10852 4446 10908
rect 4446 10852 4450 10908
rect 4386 10848 4450 10852
rect 4466 10908 4530 10912
rect 4466 10852 4470 10908
rect 4470 10852 4526 10908
rect 4526 10852 4530 10908
rect 4466 10848 4530 10852
rect 4546 10908 4610 10912
rect 4546 10852 4550 10908
rect 4550 10852 4606 10908
rect 4606 10852 4610 10908
rect 4546 10848 4610 10852
rect 4626 10908 4690 10912
rect 4626 10852 4630 10908
rect 4630 10852 4686 10908
rect 4686 10852 4690 10908
rect 4626 10848 4690 10852
rect 11256 10908 11320 10912
rect 11256 10852 11260 10908
rect 11260 10852 11316 10908
rect 11316 10852 11320 10908
rect 11256 10848 11320 10852
rect 11336 10908 11400 10912
rect 11336 10852 11340 10908
rect 11340 10852 11396 10908
rect 11396 10852 11400 10908
rect 11336 10848 11400 10852
rect 11416 10908 11480 10912
rect 11416 10852 11420 10908
rect 11420 10852 11476 10908
rect 11476 10852 11480 10908
rect 11416 10848 11480 10852
rect 11496 10908 11560 10912
rect 11496 10852 11500 10908
rect 11500 10852 11556 10908
rect 11556 10852 11560 10908
rect 11496 10848 11560 10852
rect 18125 10908 18189 10912
rect 18125 10852 18129 10908
rect 18129 10852 18185 10908
rect 18185 10852 18189 10908
rect 18125 10848 18189 10852
rect 18205 10908 18269 10912
rect 18205 10852 18209 10908
rect 18209 10852 18265 10908
rect 18265 10852 18269 10908
rect 18205 10848 18269 10852
rect 18285 10908 18349 10912
rect 18285 10852 18289 10908
rect 18289 10852 18345 10908
rect 18345 10852 18349 10908
rect 18285 10848 18349 10852
rect 18365 10908 18429 10912
rect 18365 10852 18369 10908
rect 18369 10852 18425 10908
rect 18425 10852 18429 10908
rect 18365 10848 18429 10852
rect 7821 10364 7885 10368
rect 7821 10308 7825 10364
rect 7825 10308 7881 10364
rect 7881 10308 7885 10364
rect 7821 10304 7885 10308
rect 7901 10364 7965 10368
rect 7901 10308 7905 10364
rect 7905 10308 7961 10364
rect 7961 10308 7965 10364
rect 7901 10304 7965 10308
rect 7981 10364 8045 10368
rect 7981 10308 7985 10364
rect 7985 10308 8041 10364
rect 8041 10308 8045 10364
rect 7981 10304 8045 10308
rect 8061 10364 8125 10368
rect 8061 10308 8065 10364
rect 8065 10308 8121 10364
rect 8121 10308 8125 10364
rect 8061 10304 8125 10308
rect 14690 10364 14754 10368
rect 14690 10308 14694 10364
rect 14694 10308 14750 10364
rect 14750 10308 14754 10364
rect 14690 10304 14754 10308
rect 14770 10364 14834 10368
rect 14770 10308 14774 10364
rect 14774 10308 14830 10364
rect 14830 10308 14834 10364
rect 14770 10304 14834 10308
rect 14850 10364 14914 10368
rect 14850 10308 14854 10364
rect 14854 10308 14910 10364
rect 14910 10308 14914 10364
rect 14850 10304 14914 10308
rect 14930 10364 14994 10368
rect 14930 10308 14934 10364
rect 14934 10308 14990 10364
rect 14990 10308 14994 10364
rect 14930 10304 14994 10308
rect 4386 9820 4450 9824
rect 4386 9764 4390 9820
rect 4390 9764 4446 9820
rect 4446 9764 4450 9820
rect 4386 9760 4450 9764
rect 4466 9820 4530 9824
rect 4466 9764 4470 9820
rect 4470 9764 4526 9820
rect 4526 9764 4530 9820
rect 4466 9760 4530 9764
rect 4546 9820 4610 9824
rect 4546 9764 4550 9820
rect 4550 9764 4606 9820
rect 4606 9764 4610 9820
rect 4546 9760 4610 9764
rect 4626 9820 4690 9824
rect 4626 9764 4630 9820
rect 4630 9764 4686 9820
rect 4686 9764 4690 9820
rect 4626 9760 4690 9764
rect 11256 9820 11320 9824
rect 11256 9764 11260 9820
rect 11260 9764 11316 9820
rect 11316 9764 11320 9820
rect 11256 9760 11320 9764
rect 11336 9820 11400 9824
rect 11336 9764 11340 9820
rect 11340 9764 11396 9820
rect 11396 9764 11400 9820
rect 11336 9760 11400 9764
rect 11416 9820 11480 9824
rect 11416 9764 11420 9820
rect 11420 9764 11476 9820
rect 11476 9764 11480 9820
rect 11416 9760 11480 9764
rect 11496 9820 11560 9824
rect 11496 9764 11500 9820
rect 11500 9764 11556 9820
rect 11556 9764 11560 9820
rect 11496 9760 11560 9764
rect 18125 9820 18189 9824
rect 18125 9764 18129 9820
rect 18129 9764 18185 9820
rect 18185 9764 18189 9820
rect 18125 9760 18189 9764
rect 18205 9820 18269 9824
rect 18205 9764 18209 9820
rect 18209 9764 18265 9820
rect 18265 9764 18269 9820
rect 18205 9760 18269 9764
rect 18285 9820 18349 9824
rect 18285 9764 18289 9820
rect 18289 9764 18345 9820
rect 18345 9764 18349 9820
rect 18285 9760 18349 9764
rect 18365 9820 18429 9824
rect 18365 9764 18369 9820
rect 18369 9764 18425 9820
rect 18425 9764 18429 9820
rect 18365 9760 18429 9764
rect 7821 9276 7885 9280
rect 7821 9220 7825 9276
rect 7825 9220 7881 9276
rect 7881 9220 7885 9276
rect 7821 9216 7885 9220
rect 7901 9276 7965 9280
rect 7901 9220 7905 9276
rect 7905 9220 7961 9276
rect 7961 9220 7965 9276
rect 7901 9216 7965 9220
rect 7981 9276 8045 9280
rect 7981 9220 7985 9276
rect 7985 9220 8041 9276
rect 8041 9220 8045 9276
rect 7981 9216 8045 9220
rect 8061 9276 8125 9280
rect 8061 9220 8065 9276
rect 8065 9220 8121 9276
rect 8121 9220 8125 9276
rect 8061 9216 8125 9220
rect 14690 9276 14754 9280
rect 14690 9220 14694 9276
rect 14694 9220 14750 9276
rect 14750 9220 14754 9276
rect 14690 9216 14754 9220
rect 14770 9276 14834 9280
rect 14770 9220 14774 9276
rect 14774 9220 14830 9276
rect 14830 9220 14834 9276
rect 14770 9216 14834 9220
rect 14850 9276 14914 9280
rect 14850 9220 14854 9276
rect 14854 9220 14910 9276
rect 14910 9220 14914 9276
rect 14850 9216 14914 9220
rect 14930 9276 14994 9280
rect 14930 9220 14934 9276
rect 14934 9220 14990 9276
rect 14990 9220 14994 9276
rect 14930 9216 14994 9220
rect 4386 8732 4450 8736
rect 4386 8676 4390 8732
rect 4390 8676 4446 8732
rect 4446 8676 4450 8732
rect 4386 8672 4450 8676
rect 4466 8732 4530 8736
rect 4466 8676 4470 8732
rect 4470 8676 4526 8732
rect 4526 8676 4530 8732
rect 4466 8672 4530 8676
rect 4546 8732 4610 8736
rect 4546 8676 4550 8732
rect 4550 8676 4606 8732
rect 4606 8676 4610 8732
rect 4546 8672 4610 8676
rect 4626 8732 4690 8736
rect 4626 8676 4630 8732
rect 4630 8676 4686 8732
rect 4686 8676 4690 8732
rect 4626 8672 4690 8676
rect 11256 8732 11320 8736
rect 11256 8676 11260 8732
rect 11260 8676 11316 8732
rect 11316 8676 11320 8732
rect 11256 8672 11320 8676
rect 11336 8732 11400 8736
rect 11336 8676 11340 8732
rect 11340 8676 11396 8732
rect 11396 8676 11400 8732
rect 11336 8672 11400 8676
rect 11416 8732 11480 8736
rect 11416 8676 11420 8732
rect 11420 8676 11476 8732
rect 11476 8676 11480 8732
rect 11416 8672 11480 8676
rect 11496 8732 11560 8736
rect 11496 8676 11500 8732
rect 11500 8676 11556 8732
rect 11556 8676 11560 8732
rect 11496 8672 11560 8676
rect 18125 8732 18189 8736
rect 18125 8676 18129 8732
rect 18129 8676 18185 8732
rect 18185 8676 18189 8732
rect 18125 8672 18189 8676
rect 18205 8732 18269 8736
rect 18205 8676 18209 8732
rect 18209 8676 18265 8732
rect 18265 8676 18269 8732
rect 18205 8672 18269 8676
rect 18285 8732 18349 8736
rect 18285 8676 18289 8732
rect 18289 8676 18345 8732
rect 18345 8676 18349 8732
rect 18285 8672 18349 8676
rect 18365 8732 18429 8736
rect 18365 8676 18369 8732
rect 18369 8676 18425 8732
rect 18425 8676 18429 8732
rect 18365 8672 18429 8676
rect 7821 8188 7885 8192
rect 7821 8132 7825 8188
rect 7825 8132 7881 8188
rect 7881 8132 7885 8188
rect 7821 8128 7885 8132
rect 7901 8188 7965 8192
rect 7901 8132 7905 8188
rect 7905 8132 7961 8188
rect 7961 8132 7965 8188
rect 7901 8128 7965 8132
rect 7981 8188 8045 8192
rect 7981 8132 7985 8188
rect 7985 8132 8041 8188
rect 8041 8132 8045 8188
rect 7981 8128 8045 8132
rect 8061 8188 8125 8192
rect 8061 8132 8065 8188
rect 8065 8132 8121 8188
rect 8121 8132 8125 8188
rect 8061 8128 8125 8132
rect 14690 8188 14754 8192
rect 14690 8132 14694 8188
rect 14694 8132 14750 8188
rect 14750 8132 14754 8188
rect 14690 8128 14754 8132
rect 14770 8188 14834 8192
rect 14770 8132 14774 8188
rect 14774 8132 14830 8188
rect 14830 8132 14834 8188
rect 14770 8128 14834 8132
rect 14850 8188 14914 8192
rect 14850 8132 14854 8188
rect 14854 8132 14910 8188
rect 14910 8132 14914 8188
rect 14850 8128 14914 8132
rect 14930 8188 14994 8192
rect 14930 8132 14934 8188
rect 14934 8132 14990 8188
rect 14990 8132 14994 8188
rect 14930 8128 14994 8132
rect 4386 7644 4450 7648
rect 4386 7588 4390 7644
rect 4390 7588 4446 7644
rect 4446 7588 4450 7644
rect 4386 7584 4450 7588
rect 4466 7644 4530 7648
rect 4466 7588 4470 7644
rect 4470 7588 4526 7644
rect 4526 7588 4530 7644
rect 4466 7584 4530 7588
rect 4546 7644 4610 7648
rect 4546 7588 4550 7644
rect 4550 7588 4606 7644
rect 4606 7588 4610 7644
rect 4546 7584 4610 7588
rect 4626 7644 4690 7648
rect 4626 7588 4630 7644
rect 4630 7588 4686 7644
rect 4686 7588 4690 7644
rect 4626 7584 4690 7588
rect 11256 7644 11320 7648
rect 11256 7588 11260 7644
rect 11260 7588 11316 7644
rect 11316 7588 11320 7644
rect 11256 7584 11320 7588
rect 11336 7644 11400 7648
rect 11336 7588 11340 7644
rect 11340 7588 11396 7644
rect 11396 7588 11400 7644
rect 11336 7584 11400 7588
rect 11416 7644 11480 7648
rect 11416 7588 11420 7644
rect 11420 7588 11476 7644
rect 11476 7588 11480 7644
rect 11416 7584 11480 7588
rect 11496 7644 11560 7648
rect 11496 7588 11500 7644
rect 11500 7588 11556 7644
rect 11556 7588 11560 7644
rect 11496 7584 11560 7588
rect 18125 7644 18189 7648
rect 18125 7588 18129 7644
rect 18129 7588 18185 7644
rect 18185 7588 18189 7644
rect 18125 7584 18189 7588
rect 18205 7644 18269 7648
rect 18205 7588 18209 7644
rect 18209 7588 18265 7644
rect 18265 7588 18269 7644
rect 18205 7584 18269 7588
rect 18285 7644 18349 7648
rect 18285 7588 18289 7644
rect 18289 7588 18345 7644
rect 18345 7588 18349 7644
rect 18285 7584 18349 7588
rect 18365 7644 18429 7648
rect 18365 7588 18369 7644
rect 18369 7588 18425 7644
rect 18425 7588 18429 7644
rect 18365 7584 18429 7588
rect 7821 7100 7885 7104
rect 7821 7044 7825 7100
rect 7825 7044 7881 7100
rect 7881 7044 7885 7100
rect 7821 7040 7885 7044
rect 7901 7100 7965 7104
rect 7901 7044 7905 7100
rect 7905 7044 7961 7100
rect 7961 7044 7965 7100
rect 7901 7040 7965 7044
rect 7981 7100 8045 7104
rect 7981 7044 7985 7100
rect 7985 7044 8041 7100
rect 8041 7044 8045 7100
rect 7981 7040 8045 7044
rect 8061 7100 8125 7104
rect 8061 7044 8065 7100
rect 8065 7044 8121 7100
rect 8121 7044 8125 7100
rect 8061 7040 8125 7044
rect 14690 7100 14754 7104
rect 14690 7044 14694 7100
rect 14694 7044 14750 7100
rect 14750 7044 14754 7100
rect 14690 7040 14754 7044
rect 14770 7100 14834 7104
rect 14770 7044 14774 7100
rect 14774 7044 14830 7100
rect 14830 7044 14834 7100
rect 14770 7040 14834 7044
rect 14850 7100 14914 7104
rect 14850 7044 14854 7100
rect 14854 7044 14910 7100
rect 14910 7044 14914 7100
rect 14850 7040 14914 7044
rect 14930 7100 14994 7104
rect 14930 7044 14934 7100
rect 14934 7044 14990 7100
rect 14990 7044 14994 7100
rect 14930 7040 14994 7044
rect 4386 6556 4450 6560
rect 4386 6500 4390 6556
rect 4390 6500 4446 6556
rect 4446 6500 4450 6556
rect 4386 6496 4450 6500
rect 4466 6556 4530 6560
rect 4466 6500 4470 6556
rect 4470 6500 4526 6556
rect 4526 6500 4530 6556
rect 4466 6496 4530 6500
rect 4546 6556 4610 6560
rect 4546 6500 4550 6556
rect 4550 6500 4606 6556
rect 4606 6500 4610 6556
rect 4546 6496 4610 6500
rect 4626 6556 4690 6560
rect 4626 6500 4630 6556
rect 4630 6500 4686 6556
rect 4686 6500 4690 6556
rect 4626 6496 4690 6500
rect 11256 6556 11320 6560
rect 11256 6500 11260 6556
rect 11260 6500 11316 6556
rect 11316 6500 11320 6556
rect 11256 6496 11320 6500
rect 11336 6556 11400 6560
rect 11336 6500 11340 6556
rect 11340 6500 11396 6556
rect 11396 6500 11400 6556
rect 11336 6496 11400 6500
rect 11416 6556 11480 6560
rect 11416 6500 11420 6556
rect 11420 6500 11476 6556
rect 11476 6500 11480 6556
rect 11416 6496 11480 6500
rect 11496 6556 11560 6560
rect 11496 6500 11500 6556
rect 11500 6500 11556 6556
rect 11556 6500 11560 6556
rect 11496 6496 11560 6500
rect 18125 6556 18189 6560
rect 18125 6500 18129 6556
rect 18129 6500 18185 6556
rect 18185 6500 18189 6556
rect 18125 6496 18189 6500
rect 18205 6556 18269 6560
rect 18205 6500 18209 6556
rect 18209 6500 18265 6556
rect 18265 6500 18269 6556
rect 18205 6496 18269 6500
rect 18285 6556 18349 6560
rect 18285 6500 18289 6556
rect 18289 6500 18345 6556
rect 18345 6500 18349 6556
rect 18285 6496 18349 6500
rect 18365 6556 18429 6560
rect 18365 6500 18369 6556
rect 18369 6500 18425 6556
rect 18425 6500 18429 6556
rect 18365 6496 18429 6500
rect 7821 6012 7885 6016
rect 7821 5956 7825 6012
rect 7825 5956 7881 6012
rect 7881 5956 7885 6012
rect 7821 5952 7885 5956
rect 7901 6012 7965 6016
rect 7901 5956 7905 6012
rect 7905 5956 7961 6012
rect 7961 5956 7965 6012
rect 7901 5952 7965 5956
rect 7981 6012 8045 6016
rect 7981 5956 7985 6012
rect 7985 5956 8041 6012
rect 8041 5956 8045 6012
rect 7981 5952 8045 5956
rect 8061 6012 8125 6016
rect 8061 5956 8065 6012
rect 8065 5956 8121 6012
rect 8121 5956 8125 6012
rect 8061 5952 8125 5956
rect 14690 6012 14754 6016
rect 14690 5956 14694 6012
rect 14694 5956 14750 6012
rect 14750 5956 14754 6012
rect 14690 5952 14754 5956
rect 14770 6012 14834 6016
rect 14770 5956 14774 6012
rect 14774 5956 14830 6012
rect 14830 5956 14834 6012
rect 14770 5952 14834 5956
rect 14850 6012 14914 6016
rect 14850 5956 14854 6012
rect 14854 5956 14910 6012
rect 14910 5956 14914 6012
rect 14850 5952 14914 5956
rect 14930 6012 14994 6016
rect 14930 5956 14934 6012
rect 14934 5956 14990 6012
rect 14990 5956 14994 6012
rect 14930 5952 14994 5956
rect 4386 5468 4450 5472
rect 4386 5412 4390 5468
rect 4390 5412 4446 5468
rect 4446 5412 4450 5468
rect 4386 5408 4450 5412
rect 4466 5468 4530 5472
rect 4466 5412 4470 5468
rect 4470 5412 4526 5468
rect 4526 5412 4530 5468
rect 4466 5408 4530 5412
rect 4546 5468 4610 5472
rect 4546 5412 4550 5468
rect 4550 5412 4606 5468
rect 4606 5412 4610 5468
rect 4546 5408 4610 5412
rect 4626 5468 4690 5472
rect 4626 5412 4630 5468
rect 4630 5412 4686 5468
rect 4686 5412 4690 5468
rect 4626 5408 4690 5412
rect 11256 5468 11320 5472
rect 11256 5412 11260 5468
rect 11260 5412 11316 5468
rect 11316 5412 11320 5468
rect 11256 5408 11320 5412
rect 11336 5468 11400 5472
rect 11336 5412 11340 5468
rect 11340 5412 11396 5468
rect 11396 5412 11400 5468
rect 11336 5408 11400 5412
rect 11416 5468 11480 5472
rect 11416 5412 11420 5468
rect 11420 5412 11476 5468
rect 11476 5412 11480 5468
rect 11416 5408 11480 5412
rect 11496 5468 11560 5472
rect 11496 5412 11500 5468
rect 11500 5412 11556 5468
rect 11556 5412 11560 5468
rect 11496 5408 11560 5412
rect 18125 5468 18189 5472
rect 18125 5412 18129 5468
rect 18129 5412 18185 5468
rect 18185 5412 18189 5468
rect 18125 5408 18189 5412
rect 18205 5468 18269 5472
rect 18205 5412 18209 5468
rect 18209 5412 18265 5468
rect 18265 5412 18269 5468
rect 18205 5408 18269 5412
rect 18285 5468 18349 5472
rect 18285 5412 18289 5468
rect 18289 5412 18345 5468
rect 18345 5412 18349 5468
rect 18285 5408 18349 5412
rect 18365 5468 18429 5472
rect 18365 5412 18369 5468
rect 18369 5412 18425 5468
rect 18425 5412 18429 5468
rect 18365 5408 18429 5412
rect 7821 4924 7885 4928
rect 7821 4868 7825 4924
rect 7825 4868 7881 4924
rect 7881 4868 7885 4924
rect 7821 4864 7885 4868
rect 7901 4924 7965 4928
rect 7901 4868 7905 4924
rect 7905 4868 7961 4924
rect 7961 4868 7965 4924
rect 7901 4864 7965 4868
rect 7981 4924 8045 4928
rect 7981 4868 7985 4924
rect 7985 4868 8041 4924
rect 8041 4868 8045 4924
rect 7981 4864 8045 4868
rect 8061 4924 8125 4928
rect 8061 4868 8065 4924
rect 8065 4868 8121 4924
rect 8121 4868 8125 4924
rect 8061 4864 8125 4868
rect 14690 4924 14754 4928
rect 14690 4868 14694 4924
rect 14694 4868 14750 4924
rect 14750 4868 14754 4924
rect 14690 4864 14754 4868
rect 14770 4924 14834 4928
rect 14770 4868 14774 4924
rect 14774 4868 14830 4924
rect 14830 4868 14834 4924
rect 14770 4864 14834 4868
rect 14850 4924 14914 4928
rect 14850 4868 14854 4924
rect 14854 4868 14910 4924
rect 14910 4868 14914 4924
rect 14850 4864 14914 4868
rect 14930 4924 14994 4928
rect 14930 4868 14934 4924
rect 14934 4868 14990 4924
rect 14990 4868 14994 4924
rect 14930 4864 14994 4868
rect 4386 4380 4450 4384
rect 4386 4324 4390 4380
rect 4390 4324 4446 4380
rect 4446 4324 4450 4380
rect 4386 4320 4450 4324
rect 4466 4380 4530 4384
rect 4466 4324 4470 4380
rect 4470 4324 4526 4380
rect 4526 4324 4530 4380
rect 4466 4320 4530 4324
rect 4546 4380 4610 4384
rect 4546 4324 4550 4380
rect 4550 4324 4606 4380
rect 4606 4324 4610 4380
rect 4546 4320 4610 4324
rect 4626 4380 4690 4384
rect 4626 4324 4630 4380
rect 4630 4324 4686 4380
rect 4686 4324 4690 4380
rect 4626 4320 4690 4324
rect 11256 4380 11320 4384
rect 11256 4324 11260 4380
rect 11260 4324 11316 4380
rect 11316 4324 11320 4380
rect 11256 4320 11320 4324
rect 11336 4380 11400 4384
rect 11336 4324 11340 4380
rect 11340 4324 11396 4380
rect 11396 4324 11400 4380
rect 11336 4320 11400 4324
rect 11416 4380 11480 4384
rect 11416 4324 11420 4380
rect 11420 4324 11476 4380
rect 11476 4324 11480 4380
rect 11416 4320 11480 4324
rect 11496 4380 11560 4384
rect 11496 4324 11500 4380
rect 11500 4324 11556 4380
rect 11556 4324 11560 4380
rect 11496 4320 11560 4324
rect 18125 4380 18189 4384
rect 18125 4324 18129 4380
rect 18129 4324 18185 4380
rect 18185 4324 18189 4380
rect 18125 4320 18189 4324
rect 18205 4380 18269 4384
rect 18205 4324 18209 4380
rect 18209 4324 18265 4380
rect 18265 4324 18269 4380
rect 18205 4320 18269 4324
rect 18285 4380 18349 4384
rect 18285 4324 18289 4380
rect 18289 4324 18345 4380
rect 18345 4324 18349 4380
rect 18285 4320 18349 4324
rect 18365 4380 18429 4384
rect 18365 4324 18369 4380
rect 18369 4324 18425 4380
rect 18425 4324 18429 4380
rect 18365 4320 18429 4324
rect 7821 3836 7885 3840
rect 7821 3780 7825 3836
rect 7825 3780 7881 3836
rect 7881 3780 7885 3836
rect 7821 3776 7885 3780
rect 7901 3836 7965 3840
rect 7901 3780 7905 3836
rect 7905 3780 7961 3836
rect 7961 3780 7965 3836
rect 7901 3776 7965 3780
rect 7981 3836 8045 3840
rect 7981 3780 7985 3836
rect 7985 3780 8041 3836
rect 8041 3780 8045 3836
rect 7981 3776 8045 3780
rect 8061 3836 8125 3840
rect 8061 3780 8065 3836
rect 8065 3780 8121 3836
rect 8121 3780 8125 3836
rect 8061 3776 8125 3780
rect 14690 3836 14754 3840
rect 14690 3780 14694 3836
rect 14694 3780 14750 3836
rect 14750 3780 14754 3836
rect 14690 3776 14754 3780
rect 14770 3836 14834 3840
rect 14770 3780 14774 3836
rect 14774 3780 14830 3836
rect 14830 3780 14834 3836
rect 14770 3776 14834 3780
rect 14850 3836 14914 3840
rect 14850 3780 14854 3836
rect 14854 3780 14910 3836
rect 14910 3780 14914 3836
rect 14850 3776 14914 3780
rect 14930 3836 14994 3840
rect 14930 3780 14934 3836
rect 14934 3780 14990 3836
rect 14990 3780 14994 3836
rect 14930 3776 14994 3780
rect 4386 3292 4450 3296
rect 4386 3236 4390 3292
rect 4390 3236 4446 3292
rect 4446 3236 4450 3292
rect 4386 3232 4450 3236
rect 4466 3292 4530 3296
rect 4466 3236 4470 3292
rect 4470 3236 4526 3292
rect 4526 3236 4530 3292
rect 4466 3232 4530 3236
rect 4546 3292 4610 3296
rect 4546 3236 4550 3292
rect 4550 3236 4606 3292
rect 4606 3236 4610 3292
rect 4546 3232 4610 3236
rect 4626 3292 4690 3296
rect 4626 3236 4630 3292
rect 4630 3236 4686 3292
rect 4686 3236 4690 3292
rect 4626 3232 4690 3236
rect 11256 3292 11320 3296
rect 11256 3236 11260 3292
rect 11260 3236 11316 3292
rect 11316 3236 11320 3292
rect 11256 3232 11320 3236
rect 11336 3292 11400 3296
rect 11336 3236 11340 3292
rect 11340 3236 11396 3292
rect 11396 3236 11400 3292
rect 11336 3232 11400 3236
rect 11416 3292 11480 3296
rect 11416 3236 11420 3292
rect 11420 3236 11476 3292
rect 11476 3236 11480 3292
rect 11416 3232 11480 3236
rect 11496 3292 11560 3296
rect 11496 3236 11500 3292
rect 11500 3236 11556 3292
rect 11556 3236 11560 3292
rect 11496 3232 11560 3236
rect 18125 3292 18189 3296
rect 18125 3236 18129 3292
rect 18129 3236 18185 3292
rect 18185 3236 18189 3292
rect 18125 3232 18189 3236
rect 18205 3292 18269 3296
rect 18205 3236 18209 3292
rect 18209 3236 18265 3292
rect 18265 3236 18269 3292
rect 18205 3232 18269 3236
rect 18285 3292 18349 3296
rect 18285 3236 18289 3292
rect 18289 3236 18345 3292
rect 18345 3236 18349 3292
rect 18285 3232 18349 3236
rect 18365 3292 18429 3296
rect 18365 3236 18369 3292
rect 18369 3236 18425 3292
rect 18425 3236 18429 3292
rect 18365 3232 18429 3236
rect 7821 2748 7885 2752
rect 7821 2692 7825 2748
rect 7825 2692 7881 2748
rect 7881 2692 7885 2748
rect 7821 2688 7885 2692
rect 7901 2748 7965 2752
rect 7901 2692 7905 2748
rect 7905 2692 7961 2748
rect 7961 2692 7965 2748
rect 7901 2688 7965 2692
rect 7981 2748 8045 2752
rect 7981 2692 7985 2748
rect 7985 2692 8041 2748
rect 8041 2692 8045 2748
rect 7981 2688 8045 2692
rect 8061 2748 8125 2752
rect 8061 2692 8065 2748
rect 8065 2692 8121 2748
rect 8121 2692 8125 2748
rect 8061 2688 8125 2692
rect 14690 2748 14754 2752
rect 14690 2692 14694 2748
rect 14694 2692 14750 2748
rect 14750 2692 14754 2748
rect 14690 2688 14754 2692
rect 14770 2748 14834 2752
rect 14770 2692 14774 2748
rect 14774 2692 14830 2748
rect 14830 2692 14834 2748
rect 14770 2688 14834 2692
rect 14850 2748 14914 2752
rect 14850 2692 14854 2748
rect 14854 2692 14910 2748
rect 14910 2692 14914 2748
rect 14850 2688 14914 2692
rect 14930 2748 14994 2752
rect 14930 2692 14934 2748
rect 14934 2692 14990 2748
rect 14990 2692 14994 2748
rect 14930 2688 14994 2692
rect 4386 2204 4450 2208
rect 4386 2148 4390 2204
rect 4390 2148 4446 2204
rect 4446 2148 4450 2204
rect 4386 2144 4450 2148
rect 4466 2204 4530 2208
rect 4466 2148 4470 2204
rect 4470 2148 4526 2204
rect 4526 2148 4530 2204
rect 4466 2144 4530 2148
rect 4546 2204 4610 2208
rect 4546 2148 4550 2204
rect 4550 2148 4606 2204
rect 4606 2148 4610 2204
rect 4546 2144 4610 2148
rect 4626 2204 4690 2208
rect 4626 2148 4630 2204
rect 4630 2148 4686 2204
rect 4686 2148 4690 2204
rect 4626 2144 4690 2148
rect 11256 2204 11320 2208
rect 11256 2148 11260 2204
rect 11260 2148 11316 2204
rect 11316 2148 11320 2204
rect 11256 2144 11320 2148
rect 11336 2204 11400 2208
rect 11336 2148 11340 2204
rect 11340 2148 11396 2204
rect 11396 2148 11400 2204
rect 11336 2144 11400 2148
rect 11416 2204 11480 2208
rect 11416 2148 11420 2204
rect 11420 2148 11476 2204
rect 11476 2148 11480 2204
rect 11416 2144 11480 2148
rect 11496 2204 11560 2208
rect 11496 2148 11500 2204
rect 11500 2148 11556 2204
rect 11556 2148 11560 2204
rect 11496 2144 11560 2148
rect 18125 2204 18189 2208
rect 18125 2148 18129 2204
rect 18129 2148 18185 2204
rect 18185 2148 18189 2204
rect 18125 2144 18189 2148
rect 18205 2204 18269 2208
rect 18205 2148 18209 2204
rect 18209 2148 18265 2204
rect 18265 2148 18269 2204
rect 18205 2144 18269 2148
rect 18285 2204 18349 2208
rect 18285 2148 18289 2204
rect 18289 2148 18345 2204
rect 18345 2148 18349 2204
rect 18285 2144 18349 2148
rect 18365 2204 18429 2208
rect 18365 2148 18369 2204
rect 18369 2148 18425 2204
rect 18425 2148 18429 2204
rect 18365 2144 18429 2148
<< metal4 >>
rect 4378 21792 4699 22352
rect 4378 21728 4386 21792
rect 4450 21728 4466 21792
rect 4530 21728 4546 21792
rect 4610 21728 4626 21792
rect 4690 21728 4699 21792
rect 4378 20704 4699 21728
rect 4378 20640 4386 20704
rect 4450 20640 4466 20704
rect 4530 20640 4546 20704
rect 4610 20640 4626 20704
rect 4690 20640 4699 20704
rect 4378 19616 4699 20640
rect 4378 19552 4386 19616
rect 4450 19552 4466 19616
rect 4530 19552 4546 19616
rect 4610 19552 4626 19616
rect 4690 19552 4699 19616
rect 4378 19019 4699 19552
rect 4378 18783 4420 19019
rect 4656 18783 4699 19019
rect 4378 18528 4699 18783
rect 4378 18464 4386 18528
rect 4450 18464 4466 18528
rect 4530 18464 4546 18528
rect 4610 18464 4626 18528
rect 4690 18464 4699 18528
rect 4378 17440 4699 18464
rect 4378 17376 4386 17440
rect 4450 17376 4466 17440
rect 4530 17376 4546 17440
rect 4610 17376 4626 17440
rect 4690 17376 4699 17440
rect 4378 16352 4699 17376
rect 4378 16288 4386 16352
rect 4450 16288 4466 16352
rect 4530 16288 4546 16352
rect 4610 16288 4626 16352
rect 4690 16288 4699 16352
rect 4378 15264 4699 16288
rect 4378 15200 4386 15264
rect 4450 15200 4466 15264
rect 4530 15200 4546 15264
rect 4610 15200 4626 15264
rect 4690 15200 4699 15264
rect 4378 14176 4699 15200
rect 4378 14112 4386 14176
rect 4450 14112 4466 14176
rect 4530 14112 4546 14176
rect 4610 14112 4626 14176
rect 4690 14112 4699 14176
rect 4378 13088 4699 14112
rect 4378 13024 4386 13088
rect 4450 13024 4466 13088
rect 4530 13024 4546 13088
rect 4610 13024 4626 13088
rect 4690 13024 4699 13088
rect 4378 12310 4699 13024
rect 4378 12074 4420 12310
rect 4656 12074 4699 12310
rect 4378 12000 4699 12074
rect 4378 11936 4386 12000
rect 4450 11936 4466 12000
rect 4530 11936 4546 12000
rect 4610 11936 4626 12000
rect 4690 11936 4699 12000
rect 4378 10912 4699 11936
rect 4378 10848 4386 10912
rect 4450 10848 4466 10912
rect 4530 10848 4546 10912
rect 4610 10848 4626 10912
rect 4690 10848 4699 10912
rect 4378 9824 4699 10848
rect 4378 9760 4386 9824
rect 4450 9760 4466 9824
rect 4530 9760 4546 9824
rect 4610 9760 4626 9824
rect 4690 9760 4699 9824
rect 4378 8736 4699 9760
rect 4378 8672 4386 8736
rect 4450 8672 4466 8736
rect 4530 8672 4546 8736
rect 4610 8672 4626 8736
rect 4690 8672 4699 8736
rect 4378 7648 4699 8672
rect 4378 7584 4386 7648
rect 4450 7584 4466 7648
rect 4530 7584 4546 7648
rect 4610 7584 4626 7648
rect 4690 7584 4699 7648
rect 4378 6560 4699 7584
rect 4378 6496 4386 6560
rect 4450 6496 4466 6560
rect 4530 6496 4546 6560
rect 4610 6496 4626 6560
rect 4690 6496 4699 6560
rect 4378 5600 4699 6496
rect 4378 5472 4420 5600
rect 4656 5472 4699 5600
rect 4378 5408 4386 5472
rect 4690 5408 4699 5472
rect 4378 5364 4420 5408
rect 4656 5364 4699 5408
rect 4378 4384 4699 5364
rect 4378 4320 4386 4384
rect 4450 4320 4466 4384
rect 4530 4320 4546 4384
rect 4610 4320 4626 4384
rect 4690 4320 4699 4384
rect 4378 3296 4699 4320
rect 4378 3232 4386 3296
rect 4450 3232 4466 3296
rect 4530 3232 4546 3296
rect 4610 3232 4626 3296
rect 4690 3232 4699 3296
rect 4378 2208 4699 3232
rect 4378 2144 4386 2208
rect 4450 2144 4466 2208
rect 4530 2144 4546 2208
rect 4610 2144 4626 2208
rect 4690 2144 4699 2208
rect 4378 2128 4699 2144
rect 7813 22336 8133 22352
rect 7813 22272 7821 22336
rect 7885 22272 7901 22336
rect 7965 22272 7981 22336
rect 8045 22272 8061 22336
rect 8125 22272 8133 22336
rect 7813 21248 8133 22272
rect 7813 21184 7821 21248
rect 7885 21184 7901 21248
rect 7965 21184 7981 21248
rect 8045 21184 8061 21248
rect 8125 21184 8133 21248
rect 7813 20160 8133 21184
rect 7813 20096 7821 20160
rect 7885 20096 7901 20160
rect 7965 20096 7981 20160
rect 8045 20096 8061 20160
rect 8125 20096 8133 20160
rect 7813 19072 8133 20096
rect 7813 19008 7821 19072
rect 7885 19008 7901 19072
rect 7965 19008 7981 19072
rect 8045 19008 8061 19072
rect 8125 19008 8133 19072
rect 7813 17984 8133 19008
rect 7813 17920 7821 17984
rect 7885 17920 7901 17984
rect 7965 17920 7981 17984
rect 8045 17920 8061 17984
rect 8125 17920 8133 17984
rect 7813 16896 8133 17920
rect 7813 16832 7821 16896
rect 7885 16832 7901 16896
rect 7965 16832 7981 16896
rect 8045 16832 8061 16896
rect 8125 16832 8133 16896
rect 7813 15808 8133 16832
rect 7813 15744 7821 15808
rect 7885 15744 7901 15808
rect 7965 15744 7981 15808
rect 8045 15744 8061 15808
rect 8125 15744 8133 15808
rect 7813 15664 8133 15744
rect 7813 15428 7855 15664
rect 8091 15428 8133 15664
rect 7813 14720 8133 15428
rect 7813 14656 7821 14720
rect 7885 14656 7901 14720
rect 7965 14656 7981 14720
rect 8045 14656 8061 14720
rect 8125 14656 8133 14720
rect 7813 13632 8133 14656
rect 7813 13568 7821 13632
rect 7885 13568 7901 13632
rect 7965 13568 7981 13632
rect 8045 13568 8061 13632
rect 8125 13568 8133 13632
rect 7813 12544 8133 13568
rect 7813 12480 7821 12544
rect 7885 12480 7901 12544
rect 7965 12480 7981 12544
rect 8045 12480 8061 12544
rect 8125 12480 8133 12544
rect 7813 11456 8133 12480
rect 7813 11392 7821 11456
rect 7885 11392 7901 11456
rect 7965 11392 7981 11456
rect 8045 11392 8061 11456
rect 8125 11392 8133 11456
rect 7813 10368 8133 11392
rect 7813 10304 7821 10368
rect 7885 10304 7901 10368
rect 7965 10304 7981 10368
rect 8045 10304 8061 10368
rect 8125 10304 8133 10368
rect 7813 9280 8133 10304
rect 7813 9216 7821 9280
rect 7885 9216 7901 9280
rect 7965 9216 7981 9280
rect 8045 9216 8061 9280
rect 8125 9216 8133 9280
rect 7813 8955 8133 9216
rect 7813 8719 7855 8955
rect 8091 8719 8133 8955
rect 7813 8192 8133 8719
rect 7813 8128 7821 8192
rect 7885 8128 7901 8192
rect 7965 8128 7981 8192
rect 8045 8128 8061 8192
rect 8125 8128 8133 8192
rect 7813 7104 8133 8128
rect 7813 7040 7821 7104
rect 7885 7040 7901 7104
rect 7965 7040 7981 7104
rect 8045 7040 8061 7104
rect 8125 7040 8133 7104
rect 7813 6016 8133 7040
rect 7813 5952 7821 6016
rect 7885 5952 7901 6016
rect 7965 5952 7981 6016
rect 8045 5952 8061 6016
rect 8125 5952 8133 6016
rect 7813 4928 8133 5952
rect 7813 4864 7821 4928
rect 7885 4864 7901 4928
rect 7965 4864 7981 4928
rect 8045 4864 8061 4928
rect 8125 4864 8133 4928
rect 7813 3840 8133 4864
rect 7813 3776 7821 3840
rect 7885 3776 7901 3840
rect 7965 3776 7981 3840
rect 8045 3776 8061 3840
rect 8125 3776 8133 3840
rect 7813 2752 8133 3776
rect 7813 2688 7821 2752
rect 7885 2688 7901 2752
rect 7965 2688 7981 2752
rect 8045 2688 8061 2752
rect 8125 2688 8133 2752
rect 7813 2128 8133 2688
rect 11248 21792 11568 22352
rect 11248 21728 11256 21792
rect 11320 21728 11336 21792
rect 11400 21728 11416 21792
rect 11480 21728 11496 21792
rect 11560 21728 11568 21792
rect 11248 20704 11568 21728
rect 11248 20640 11256 20704
rect 11320 20640 11336 20704
rect 11400 20640 11416 20704
rect 11480 20640 11496 20704
rect 11560 20640 11568 20704
rect 11248 19616 11568 20640
rect 11248 19552 11256 19616
rect 11320 19552 11336 19616
rect 11400 19552 11416 19616
rect 11480 19552 11496 19616
rect 11560 19552 11568 19616
rect 11248 19019 11568 19552
rect 11248 18783 11290 19019
rect 11526 18783 11568 19019
rect 11248 18528 11568 18783
rect 11248 18464 11256 18528
rect 11320 18464 11336 18528
rect 11400 18464 11416 18528
rect 11480 18464 11496 18528
rect 11560 18464 11568 18528
rect 11248 17440 11568 18464
rect 11248 17376 11256 17440
rect 11320 17376 11336 17440
rect 11400 17376 11416 17440
rect 11480 17376 11496 17440
rect 11560 17376 11568 17440
rect 11248 16352 11568 17376
rect 11248 16288 11256 16352
rect 11320 16288 11336 16352
rect 11400 16288 11416 16352
rect 11480 16288 11496 16352
rect 11560 16288 11568 16352
rect 11248 15264 11568 16288
rect 11248 15200 11256 15264
rect 11320 15200 11336 15264
rect 11400 15200 11416 15264
rect 11480 15200 11496 15264
rect 11560 15200 11568 15264
rect 11248 14176 11568 15200
rect 11248 14112 11256 14176
rect 11320 14112 11336 14176
rect 11400 14112 11416 14176
rect 11480 14112 11496 14176
rect 11560 14112 11568 14176
rect 11248 13088 11568 14112
rect 11248 13024 11256 13088
rect 11320 13024 11336 13088
rect 11400 13024 11416 13088
rect 11480 13024 11496 13088
rect 11560 13024 11568 13088
rect 11248 12310 11568 13024
rect 11248 12074 11290 12310
rect 11526 12074 11568 12310
rect 11248 12000 11568 12074
rect 11248 11936 11256 12000
rect 11320 11936 11336 12000
rect 11400 11936 11416 12000
rect 11480 11936 11496 12000
rect 11560 11936 11568 12000
rect 11248 10912 11568 11936
rect 11248 10848 11256 10912
rect 11320 10848 11336 10912
rect 11400 10848 11416 10912
rect 11480 10848 11496 10912
rect 11560 10848 11568 10912
rect 11248 9824 11568 10848
rect 11248 9760 11256 9824
rect 11320 9760 11336 9824
rect 11400 9760 11416 9824
rect 11480 9760 11496 9824
rect 11560 9760 11568 9824
rect 11248 8736 11568 9760
rect 11248 8672 11256 8736
rect 11320 8672 11336 8736
rect 11400 8672 11416 8736
rect 11480 8672 11496 8736
rect 11560 8672 11568 8736
rect 11248 7648 11568 8672
rect 11248 7584 11256 7648
rect 11320 7584 11336 7648
rect 11400 7584 11416 7648
rect 11480 7584 11496 7648
rect 11560 7584 11568 7648
rect 11248 6560 11568 7584
rect 11248 6496 11256 6560
rect 11320 6496 11336 6560
rect 11400 6496 11416 6560
rect 11480 6496 11496 6560
rect 11560 6496 11568 6560
rect 11248 5600 11568 6496
rect 11248 5472 11290 5600
rect 11526 5472 11568 5600
rect 11248 5408 11256 5472
rect 11560 5408 11568 5472
rect 11248 5364 11290 5408
rect 11526 5364 11568 5408
rect 11248 4384 11568 5364
rect 11248 4320 11256 4384
rect 11320 4320 11336 4384
rect 11400 4320 11416 4384
rect 11480 4320 11496 4384
rect 11560 4320 11568 4384
rect 11248 3296 11568 4320
rect 11248 3232 11256 3296
rect 11320 3232 11336 3296
rect 11400 3232 11416 3296
rect 11480 3232 11496 3296
rect 11560 3232 11568 3296
rect 11248 2208 11568 3232
rect 11248 2144 11256 2208
rect 11320 2144 11336 2208
rect 11400 2144 11416 2208
rect 11480 2144 11496 2208
rect 11560 2144 11568 2208
rect 11248 2128 11568 2144
rect 14682 22336 15003 22352
rect 14682 22272 14690 22336
rect 14754 22272 14770 22336
rect 14834 22272 14850 22336
rect 14914 22272 14930 22336
rect 14994 22272 15003 22336
rect 14682 21248 15003 22272
rect 14682 21184 14690 21248
rect 14754 21184 14770 21248
rect 14834 21184 14850 21248
rect 14914 21184 14930 21248
rect 14994 21184 15003 21248
rect 14682 20160 15003 21184
rect 14682 20096 14690 20160
rect 14754 20096 14770 20160
rect 14834 20096 14850 20160
rect 14914 20096 14930 20160
rect 14994 20096 15003 20160
rect 14682 19072 15003 20096
rect 14682 19008 14690 19072
rect 14754 19008 14770 19072
rect 14834 19008 14850 19072
rect 14914 19008 14930 19072
rect 14994 19008 15003 19072
rect 14682 17984 15003 19008
rect 14682 17920 14690 17984
rect 14754 17920 14770 17984
rect 14834 17920 14850 17984
rect 14914 17920 14930 17984
rect 14994 17920 15003 17984
rect 14682 16896 15003 17920
rect 14682 16832 14690 16896
rect 14754 16832 14770 16896
rect 14834 16832 14850 16896
rect 14914 16832 14930 16896
rect 14994 16832 15003 16896
rect 14682 15808 15003 16832
rect 14682 15744 14690 15808
rect 14754 15744 14770 15808
rect 14834 15744 14850 15808
rect 14914 15744 14930 15808
rect 14994 15744 15003 15808
rect 14682 15664 15003 15744
rect 14682 15428 14724 15664
rect 14960 15428 15003 15664
rect 14682 14720 15003 15428
rect 14682 14656 14690 14720
rect 14754 14656 14770 14720
rect 14834 14656 14850 14720
rect 14914 14656 14930 14720
rect 14994 14656 15003 14720
rect 14682 13632 15003 14656
rect 14682 13568 14690 13632
rect 14754 13568 14770 13632
rect 14834 13568 14850 13632
rect 14914 13568 14930 13632
rect 14994 13568 15003 13632
rect 14682 12544 15003 13568
rect 14682 12480 14690 12544
rect 14754 12480 14770 12544
rect 14834 12480 14850 12544
rect 14914 12480 14930 12544
rect 14994 12480 15003 12544
rect 14682 11456 15003 12480
rect 14682 11392 14690 11456
rect 14754 11392 14770 11456
rect 14834 11392 14850 11456
rect 14914 11392 14930 11456
rect 14994 11392 15003 11456
rect 14682 10368 15003 11392
rect 14682 10304 14690 10368
rect 14754 10304 14770 10368
rect 14834 10304 14850 10368
rect 14914 10304 14930 10368
rect 14994 10304 15003 10368
rect 14682 9280 15003 10304
rect 14682 9216 14690 9280
rect 14754 9216 14770 9280
rect 14834 9216 14850 9280
rect 14914 9216 14930 9280
rect 14994 9216 15003 9280
rect 14682 8955 15003 9216
rect 14682 8719 14724 8955
rect 14960 8719 15003 8955
rect 14682 8192 15003 8719
rect 14682 8128 14690 8192
rect 14754 8128 14770 8192
rect 14834 8128 14850 8192
rect 14914 8128 14930 8192
rect 14994 8128 15003 8192
rect 14682 7104 15003 8128
rect 14682 7040 14690 7104
rect 14754 7040 14770 7104
rect 14834 7040 14850 7104
rect 14914 7040 14930 7104
rect 14994 7040 15003 7104
rect 14682 6016 15003 7040
rect 14682 5952 14690 6016
rect 14754 5952 14770 6016
rect 14834 5952 14850 6016
rect 14914 5952 14930 6016
rect 14994 5952 15003 6016
rect 14682 4928 15003 5952
rect 14682 4864 14690 4928
rect 14754 4864 14770 4928
rect 14834 4864 14850 4928
rect 14914 4864 14930 4928
rect 14994 4864 15003 4928
rect 14682 3840 15003 4864
rect 14682 3776 14690 3840
rect 14754 3776 14770 3840
rect 14834 3776 14850 3840
rect 14914 3776 14930 3840
rect 14994 3776 15003 3840
rect 14682 2752 15003 3776
rect 14682 2688 14690 2752
rect 14754 2688 14770 2752
rect 14834 2688 14850 2752
rect 14914 2688 14930 2752
rect 14994 2688 15003 2752
rect 14682 2128 15003 2688
rect 18117 21792 18437 22352
rect 18117 21728 18125 21792
rect 18189 21728 18205 21792
rect 18269 21728 18285 21792
rect 18349 21728 18365 21792
rect 18429 21728 18437 21792
rect 18117 20704 18437 21728
rect 18117 20640 18125 20704
rect 18189 20640 18205 20704
rect 18269 20640 18285 20704
rect 18349 20640 18365 20704
rect 18429 20640 18437 20704
rect 18117 19616 18437 20640
rect 18117 19552 18125 19616
rect 18189 19552 18205 19616
rect 18269 19552 18285 19616
rect 18349 19552 18365 19616
rect 18429 19552 18437 19616
rect 18117 19019 18437 19552
rect 18117 18783 18159 19019
rect 18395 18783 18437 19019
rect 18117 18528 18437 18783
rect 18117 18464 18125 18528
rect 18189 18464 18205 18528
rect 18269 18464 18285 18528
rect 18349 18464 18365 18528
rect 18429 18464 18437 18528
rect 18117 17440 18437 18464
rect 18117 17376 18125 17440
rect 18189 17376 18205 17440
rect 18269 17376 18285 17440
rect 18349 17376 18365 17440
rect 18429 17376 18437 17440
rect 18117 16352 18437 17376
rect 18117 16288 18125 16352
rect 18189 16288 18205 16352
rect 18269 16288 18285 16352
rect 18349 16288 18365 16352
rect 18429 16288 18437 16352
rect 18117 15264 18437 16288
rect 18117 15200 18125 15264
rect 18189 15200 18205 15264
rect 18269 15200 18285 15264
rect 18349 15200 18365 15264
rect 18429 15200 18437 15264
rect 18117 14176 18437 15200
rect 18117 14112 18125 14176
rect 18189 14112 18205 14176
rect 18269 14112 18285 14176
rect 18349 14112 18365 14176
rect 18429 14112 18437 14176
rect 18117 13088 18437 14112
rect 18117 13024 18125 13088
rect 18189 13024 18205 13088
rect 18269 13024 18285 13088
rect 18349 13024 18365 13088
rect 18429 13024 18437 13088
rect 18117 12310 18437 13024
rect 18117 12074 18159 12310
rect 18395 12074 18437 12310
rect 18117 12000 18437 12074
rect 18117 11936 18125 12000
rect 18189 11936 18205 12000
rect 18269 11936 18285 12000
rect 18349 11936 18365 12000
rect 18429 11936 18437 12000
rect 18117 10912 18437 11936
rect 18117 10848 18125 10912
rect 18189 10848 18205 10912
rect 18269 10848 18285 10912
rect 18349 10848 18365 10912
rect 18429 10848 18437 10912
rect 18117 9824 18437 10848
rect 18117 9760 18125 9824
rect 18189 9760 18205 9824
rect 18269 9760 18285 9824
rect 18349 9760 18365 9824
rect 18429 9760 18437 9824
rect 18117 8736 18437 9760
rect 18117 8672 18125 8736
rect 18189 8672 18205 8736
rect 18269 8672 18285 8736
rect 18349 8672 18365 8736
rect 18429 8672 18437 8736
rect 18117 7648 18437 8672
rect 18117 7584 18125 7648
rect 18189 7584 18205 7648
rect 18269 7584 18285 7648
rect 18349 7584 18365 7648
rect 18429 7584 18437 7648
rect 18117 6560 18437 7584
rect 18117 6496 18125 6560
rect 18189 6496 18205 6560
rect 18269 6496 18285 6560
rect 18349 6496 18365 6560
rect 18429 6496 18437 6560
rect 18117 5600 18437 6496
rect 18117 5472 18159 5600
rect 18395 5472 18437 5600
rect 18117 5408 18125 5472
rect 18429 5408 18437 5472
rect 18117 5364 18159 5408
rect 18395 5364 18437 5408
rect 18117 4384 18437 5364
rect 18117 4320 18125 4384
rect 18189 4320 18205 4384
rect 18269 4320 18285 4384
rect 18349 4320 18365 4384
rect 18429 4320 18437 4384
rect 18117 3296 18437 4320
rect 18117 3232 18125 3296
rect 18189 3232 18205 3296
rect 18269 3232 18285 3296
rect 18349 3232 18365 3296
rect 18429 3232 18437 3296
rect 18117 2208 18437 3232
rect 18117 2144 18125 2208
rect 18189 2144 18205 2208
rect 18269 2144 18285 2208
rect 18349 2144 18365 2208
rect 18429 2144 18437 2208
rect 18117 2128 18437 2144
<< via4 >>
rect 4420 18783 4656 19019
rect 4420 12074 4656 12310
rect 4420 5472 4656 5600
rect 4420 5408 4450 5472
rect 4450 5408 4466 5472
rect 4466 5408 4530 5472
rect 4530 5408 4546 5472
rect 4546 5408 4610 5472
rect 4610 5408 4626 5472
rect 4626 5408 4656 5472
rect 4420 5364 4656 5408
rect 7855 15428 8091 15664
rect 7855 8719 8091 8955
rect 11290 18783 11526 19019
rect 11290 12074 11526 12310
rect 11290 5472 11526 5600
rect 11290 5408 11320 5472
rect 11320 5408 11336 5472
rect 11336 5408 11400 5472
rect 11400 5408 11416 5472
rect 11416 5408 11480 5472
rect 11480 5408 11496 5472
rect 11496 5408 11526 5472
rect 11290 5364 11526 5408
rect 14724 15428 14960 15664
rect 14724 8719 14960 8955
rect 18159 18783 18395 19019
rect 18159 12074 18395 12310
rect 18159 5472 18395 5600
rect 18159 5408 18189 5472
rect 18189 5408 18205 5472
rect 18205 5408 18269 5472
rect 18269 5408 18285 5472
rect 18285 5408 18349 5472
rect 18349 5408 18365 5472
rect 18365 5408 18395 5472
rect 18159 5364 18395 5408
<< metal5 >>
rect 1104 19019 21712 19061
rect 1104 18783 4420 19019
rect 4656 18783 11290 19019
rect 11526 18783 18159 19019
rect 18395 18783 21712 19019
rect 1104 18741 21712 18783
rect 1104 15664 21712 15707
rect 1104 15428 7855 15664
rect 8091 15428 14724 15664
rect 14960 15428 21712 15664
rect 1104 15386 21712 15428
rect 1104 12310 21712 12352
rect 1104 12074 4420 12310
rect 4656 12074 11290 12310
rect 11526 12074 18159 12310
rect 18395 12074 21712 12310
rect 1104 12032 21712 12074
rect 1104 8955 21712 8997
rect 1104 8719 7855 8955
rect 8091 8719 14724 8955
rect 14960 8719 21712 8955
rect 1104 8677 21712 8719
rect 1104 5600 21712 5643
rect 1104 5364 4420 5600
rect 4656 5364 11290 5600
rect 11526 5364 18159 5600
rect 18395 5364 21712 5600
rect 1104 5322 21712 5364
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1614532237
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1614532237
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1614532237
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1614532237
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1614532237
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1614532237
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1614532237
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1614532237
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1614532237
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1614532237
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1614532237
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1614532237
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1614532237
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1614532237
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51
timestamp 1614532237
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1614532237
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1614532237
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1614532237
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1614532237
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1614532237
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1614532237
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1614532237
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1614532237
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1614532237
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1614532237
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1614532237
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1614532237
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1614532237
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1614532237
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1614532237
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1614532237
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1614532237
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1614532237
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1614532237
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1614532237
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1614532237
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1614532237
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1614532237
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1614532237
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1614532237
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1614532237
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1614532237
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1614532237
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1614532237
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1614532237
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1614532237
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1614532237
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1614532237
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1614532237
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1614532237
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_218
timestamp 1614532237
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1614532237
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1614532237
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_220
timestamp 1614532237
transform 1 0 21344 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1614532237
transform -1 0 21712 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1614532237
transform -1 0 21712 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1614532237
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1614532237
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1614532237
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1614532237
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1614532237
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1614532237
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1614532237
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1614532237
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1614532237
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1614532237
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1614532237
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1614532237
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1614532237
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1614532237
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1614532237
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1614532237
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1614532237
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1614532237
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1614532237
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1614532237
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1614532237
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1614532237
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_215
timestamp 1614532237
transform 1 0 20884 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1614532237
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1614532237
transform -1 0 21712 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1614532237
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1614532237
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1614532237
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1614532237
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1614532237
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1614532237
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1614532237
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1614532237
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1614532237
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1614532237
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1614532237
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1614532237
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1614532237
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1614532237
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1614532237
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1614532237
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1614532237
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1614532237
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1614532237
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1614532237
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1614532237
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1614532237
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1614532237
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_220
timestamp 1614532237
transform 1 0 21344 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1614532237
transform -1 0 21712 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1614532237
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1614532237
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1614532237
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1614532237
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1614532237
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1614532237
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1614532237
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1614532237
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1614532237
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1614532237
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1614532237
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1614532237
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1614532237
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1614532237
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1614532237
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1614532237
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1614532237
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1614532237
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1614532237
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1614532237
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1614532237
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1614532237
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_215
timestamp 1614532237
transform 1 0 20884 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1614532237
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1614532237
transform -1 0 21712 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1614532237
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1614532237
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1614532237
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1614532237
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1614532237
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1614532237
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1614532237
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1614532237
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1614532237
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1614532237
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1614532237
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1614532237
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1614532237
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1614532237
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1614532237
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1614532237
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1614532237
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1614532237
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1614532237
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1614532237
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1614532237
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1614532237
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1614532237
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_220
timestamp 1614532237
transform 1 0 21344 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1614532237
transform -1 0 21712 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1614532237
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1614532237
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1614532237
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1614532237
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1614532237
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1614532237
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1614532237
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1614532237
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1614532237
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1614532237
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1614532237
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1614532237
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1614532237
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1614532237
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1614532237
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1614532237
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1614532237
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1614532237
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1614532237
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1614532237
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1614532237
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1614532237
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1614532237
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1614532237
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1614532237
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1614532237
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1614532237
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1614532237
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1614532237
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1614532237
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1614532237
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1614532237
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1614532237
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1614532237
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1614532237
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1614532237
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1614532237
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1614532237
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1614532237
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1614532237
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1614532237
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1614532237
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1614532237
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1614532237
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1614532237
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_215
timestamp 1614532237
transform 1 0 20884 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1614532237
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_220
timestamp 1614532237
transform 1 0 21344 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1614532237
transform -1 0 21712 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1614532237
transform -1 0 21712 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1614532237
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1614532237
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1614532237
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1614532237
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1614532237
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1614532237
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1614532237
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1614532237
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1614532237
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1614532237
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1614532237
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1614532237
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1614532237
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1614532237
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1614532237
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1614532237
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1614532237
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1614532237
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1614532237
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1614532237
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1614532237
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1614532237
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_215
timestamp 1614532237
transform 1 0 20884 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1614532237
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1614532237
transform -1 0 21712 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1614532237
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1614532237
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1614532237
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1614532237
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1614532237
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1614532237
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1614532237
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1614532237
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1614532237
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1614532237
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1614532237
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1614532237
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1614532237
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1614532237
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1614532237
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1614532237
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1614532237
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1614532237
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1614532237
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1614532237
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1614532237
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1614532237
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1614532237
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_220
timestamp 1614532237
transform 1 0 21344 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1614532237
transform -1 0 21712 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1614532237
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1614532237
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1614532237
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1614532237
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1614532237
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1614532237
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1614532237
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1614532237
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1614532237
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1614532237
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1614532237
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1614532237
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1614532237
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1614532237
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1614532237
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1614532237
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1614532237
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1614532237
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1614532237
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1614532237
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1614532237
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1614532237
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_215
timestamp 1614532237
transform 1 0 20884 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1614532237
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1614532237
transform -1 0 21712 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1614532237
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1614532237
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1614532237
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1614532237
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1614532237
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1614532237
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1614532237
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1614532237
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1614532237
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1614532237
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1614532237
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1614532237
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_114
timestamp 1614532237
transform 1 0 11592 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_0
timestamp 1614532237
transform 1 0 11224 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1614532237
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1614532237
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1614532237
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1614532237
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1614532237
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1614532237
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1614532237
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1614532237
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_196
timestamp 1614532237
transform 1 0 19136 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _25_
timestamp 1614532237
transform 1 0 19228 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_213
timestamp 1614532237
transform 1 0 20700 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1614532237
transform -1 0 21712 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1614532237
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1614532237
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1614532237
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1614532237
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1614532237
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1614532237
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1614532237
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1614532237
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1614532237
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1614532237
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1614532237
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1614532237
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1614532237
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _44_
timestamp 1614532237
transform 1 0 10580 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_119
timestamp 1614532237
transform 1 0 12052 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _43_
timestamp 1614532237
transform 1 0 12788 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1614532237
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1614532237
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1614532237
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1614532237
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1614532237
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_198
timestamp 1614532237
transform 1 0 19320 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_190
timestamp 1614532237
transform 1 0 18584 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _34_
timestamp 1614532237
transform 1 0 19412 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_12_215
timestamp 1614532237
transform 1 0 20884 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_206
timestamp 1614532237
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1614532237
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1614532237
transform -1 0 21712 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1614532237
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1614532237
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1614532237
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1614532237
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1614532237
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1614532237
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1614532237
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1614532237
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1614532237
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1614532237
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1614532237
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1614532237
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1614532237
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1614532237
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1614532237
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1614532237
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1614532237
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1614532237
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1614532237
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1614532237
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1614532237
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_92
timestamp 1614532237
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_86
timestamp 1614532237
transform 1 0 9016 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1614532237
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _46_
timestamp 1614532237
transform 1 0 10028 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _41_
timestamp 1614532237
transform 1 0 9660 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_112
timestamp 1614532237
transform 1 0 11408 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_104
timestamp 1614532237
transform 1 0 10672 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_109
timestamp 1614532237
transform 1 0 11132 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _37_
timestamp 1614532237
transform 1 0 11500 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 1614532237
transform 1 0 12972 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_130
timestamp 1614532237
transform 1 0 13064 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1614532237
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1614532237
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _42_
timestamp 1614532237
transform 1 0 12420 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1614532237
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_137
timestamp 1614532237
transform 1 0 13708 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _49_
timestamp 1614532237
transform 1 0 13800 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_4  _45_
timestamp 1614532237
transform 1 0 13800 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_13_166
timestamp 1614532237
transform 1 0 16376 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_154
timestamp 1614532237
transform 1 0 15272 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1614532237
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _50_
timestamp 1614532237
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_14_184
timestamp 1614532237
transform 1 0 18032 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_178
timestamp 1614532237
transform 1 0 17480 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_170
timestamp 1614532237
transform 1 0 16744 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1614532237
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1614532237
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1614532237
transform 1 0 17480 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_6
timestamp 1614532237
transform 1 0 17664 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1614532237
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_196
timestamp 1614532237
transform 1 0 19136 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _35_
timestamp 1614532237
transform 1 0 18768 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__a2bb2o_4  _32_
timestamp 1614532237
transform 1 0 19228 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_14_215
timestamp 1614532237
transform 1 0 20884 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_206
timestamp 1614532237
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_213
timestamp 1614532237
transform 1 0 20700 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1614532237
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1614532237
transform -1 0 21712 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1614532237
transform -1 0 21712 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1614532237
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1614532237
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1614532237
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1614532237
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1614532237
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1614532237
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1614532237
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1614532237
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1614532237
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1614532237
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_86
timestamp 1614532237
transform 1 0 9016 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _47_
timestamp 1614532237
transform 1 0 9752 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_15_108
timestamp 1614532237
transform 1 0 11040 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1614532237
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1614532237
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1614532237
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _40_
timestamp 1614532237
transform 1 0 12604 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_141
timestamp 1614532237
transform 1 0 14076 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _48_
timestamp 1614532237
transform 1 0 14812 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_15_163
timestamp 1614532237
transform 1 0 16100 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_184
timestamp 1614532237
transform 1 0 18032 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_175
timestamp 1614532237
transform 1 0 17204 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_4
timestamp 1614532237
transform 1 0 18124 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1614532237
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_189
timestamp 1614532237
transform 1 0 18492 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _36_
timestamp 1614532237
transform 1 0 19228 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_213
timestamp 1614532237
transform 1 0 20700 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1614532237
transform -1 0 21712 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1614532237
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1614532237
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1614532237
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1614532237
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1614532237
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1614532237
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1614532237
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1614532237
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1614532237
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1614532237
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1614532237
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1614532237
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1614532237
transform 1 0 11132 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_1
timestamp 1614532237
transform 1 0 10764 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_126
timestamp 1614532237
transform 1 0 12696 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_121
timestamp 1614532237
transform 1 0 12236 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_3
timestamp 1614532237
transform 1 0 12328 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_2
timestamp 1614532237
transform 1 0 13432 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1614532237
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_138
timestamp 1614532237
transform 1 0 13800 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1614532237
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1614532237
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_23
timestamp 1614532237
transform 1 0 16560 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1614532237
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_184
timestamp 1614532237
transform 1 0 18032 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_172
timestamp 1614532237
transform 1 0 16928 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_15
timestamp 1614532237
transform 1 0 17664 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _39_
timestamp 1614532237
transform 1 0 18768 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_16_215
timestamp 1614532237
transform 1 0 20884 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1614532237
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1614532237
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1614532237
transform -1 0 21712 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1614532237
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1614532237
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1614532237
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1614532237
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1614532237
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1614532237
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1614532237
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1614532237
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1614532237
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1614532237
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1614532237
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1614532237
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1614532237
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1614532237
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1614532237
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1614532237
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1614532237
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1614532237
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1614532237
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1614532237
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_11
timestamp 1614532237
transform 1 0 18124 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1614532237
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_189
timestamp 1614532237
transform 1 0 18492 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _33_
timestamp 1614532237
transform 1 0 19228 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_213
timestamp 1614532237
transform 1 0 20700 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1614532237
transform -1 0 21712 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1614532237
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1614532237
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1614532237
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1614532237
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1614532237
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1614532237
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1614532237
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1614532237
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1614532237
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1614532237
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1614532237
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1614532237
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1614532237
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1614532237
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1614532237
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1614532237
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1614532237
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1614532237
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1614532237
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_178
timestamp 1614532237
transform 1 0 17480 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_191
timestamp 1614532237
transform 1 0 18676 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_186
timestamp 1614532237
transform 1 0 18216 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_19
timestamp 1614532237
transform 1 0 18308 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _38_
timestamp 1614532237
transform 1 0 19412 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_18_215
timestamp 1614532237
transform 1 0 20884 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_206
timestamp 1614532237
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1614532237
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1614532237
transform -1 0 21712 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1614532237
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1614532237
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1614532237
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1614532237
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1614532237
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1614532237
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1614532237
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1614532237
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1614532237
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1614532237
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1614532237
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1614532237
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1614532237
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1614532237
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1614532237
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1614532237
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1614532237
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1614532237
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1614532237
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1614532237
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1614532237
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1614532237
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1614532237
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1614532237
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1614532237
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1614532237
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1614532237
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1614532237
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1614532237
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1614532237
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1614532237
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1614532237
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1614532237
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1614532237
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1614532237
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1614532237
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1614532237
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1614532237
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1614532237
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1614532237
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1614532237
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1614532237
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1614532237
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_196
timestamp 1614532237
transform 1 0 19136 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_5
timestamp 1614532237
transform 1 0 19688 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_215
timestamp 1614532237
transform 1 0 20884 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_218
timestamp 1614532237
transform 1 0 21160 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_206
timestamp 1614532237
transform 1 0 20056 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1614532237
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1614532237
transform -1 0 21712 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1614532237
transform -1 0 21712 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1614532237
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1614532237
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1614532237
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1614532237
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1614532237
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1614532237
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1614532237
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1614532237
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1614532237
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1614532237
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1614532237
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1614532237
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1614532237
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1614532237
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1614532237
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1614532237
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1614532237
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1614532237
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1614532237
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1614532237
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1614532237
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1614532237
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1614532237
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_220
timestamp 1614532237
transform 1 0 21344 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1614532237
transform -1 0 21712 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1614532237
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1614532237
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1614532237
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1614532237
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1614532237
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1614532237
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1614532237
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1614532237
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1614532237
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1614532237
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1614532237
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1614532237
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1614532237
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1614532237
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1614532237
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1614532237
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1614532237
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1614532237
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1614532237
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1614532237
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1614532237
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1614532237
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_215
timestamp 1614532237
transform 1 0 20884 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1614532237
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1614532237
transform -1 0 21712 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1614532237
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1614532237
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1614532237
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1614532237
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1614532237
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1614532237
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1614532237
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1614532237
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1614532237
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1614532237
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1614532237
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1614532237
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1614532237
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1614532237
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1614532237
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1614532237
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1614532237
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1614532237
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1614532237
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1614532237
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1614532237
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1614532237
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1614532237
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_220
timestamp 1614532237
transform 1 0 21344 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1614532237
transform -1 0 21712 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1614532237
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1614532237
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1614532237
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1614532237
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1614532237
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1614532237
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1614532237
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1614532237
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1614532237
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1614532237
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1614532237
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1614532237
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1614532237
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1614532237
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1614532237
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1614532237
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1614532237
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1614532237
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1614532237
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1614532237
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1614532237
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1614532237
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_215
timestamp 1614532237
transform 1 0 20884 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1614532237
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1614532237
transform -1 0 21712 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1614532237
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1614532237
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1614532237
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1614532237
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1614532237
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1614532237
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1614532237
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1614532237
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1614532237
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1614532237
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1614532237
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1614532237
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1614532237
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1614532237
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1614532237
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1614532237
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1614532237
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1614532237
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1614532237
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1614532237
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1614532237
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1614532237
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1614532237
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_220
timestamp 1614532237
transform 1 0 21344 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1614532237
transform -1 0 21712 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_9
timestamp 1614532237
transform 1 0 1932 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1614532237
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_15
timestamp 1614532237
transform 1 0 2484 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1614532237
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1614532237
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1614532237
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _52_
timestamp 1614532237
transform 1 0 1656 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_33
timestamp 1614532237
transform 1 0 4140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_21
timestamp 1614532237
transform 1 0 3036 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1614532237
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1614532237
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_34
timestamp 1614532237
transform 1 0 3772 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_32
timestamp 1614532237
transform 1 0 2852 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_18
timestamp 1614532237
transform 1 0 2668 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1614532237
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_45
timestamp 1614532237
transform 1 0 5244 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1614532237
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1614532237
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1614532237
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1614532237
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1614532237
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1614532237
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1614532237
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1614532237
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1614532237
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1614532237
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1614532237
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1614532237
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1614532237
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1614532237
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1614532237
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1614532237
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1614532237
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1614532237
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1614532237
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1614532237
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1614532237
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1614532237
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1614532237
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1614532237
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1614532237
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1614532237
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1614532237
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1614532237
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1614532237
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1614532237
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1614532237
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1614532237
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1614532237
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_215
timestamp 1614532237
transform 1 0 20884 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1614532237
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_220
timestamp 1614532237
transform 1 0 21344 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1614532237
transform -1 0 21712 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1614532237
transform -1 0 21712 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_7
timestamp 1614532237
transform 1 0 1748 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_35
timestamp 1614532237
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1614532237
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _28_
timestamp 1614532237
transform 1 0 2484 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1614532237
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_22
timestamp 1614532237
transform 1 0 3128 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_22
timestamp 1614532237
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1614532237
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_48
timestamp 1614532237
transform 1 0 5520 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_36
timestamp 1614532237
transform 1 0 4416 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_60
timestamp 1614532237
transform 1 0 6624 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1614532237
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_72
timestamp 1614532237
transform 1 0 7728 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1614532237
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1614532237
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1614532237
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1614532237
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1614532237
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1614532237
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1614532237
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1614532237
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1614532237
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1614532237
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1614532237
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1614532237
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_215
timestamp 1614532237
transform 1 0 20884 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1614532237
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1614532237
transform -1 0 21712 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1614532237
transform 1 0 1748 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1614532237
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1614532237
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _29_
timestamp 1614532237
transform 1 0 1840 0 1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_29_22
timestamp 1614532237
transform 1 0 3128 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _53_
timestamp 1614532237
transform 1 0 3864 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_42
timestamp 1614532237
transform 1 0 4968 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1614532237
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_60
timestamp 1614532237
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_54
timestamp 1614532237
transform 1 0 6072 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1614532237
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1614532237
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1614532237
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1614532237
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1614532237
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1614532237
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1614532237
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1614532237
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1614532237
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1614532237
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1614532237
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1614532237
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1614532237
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1614532237
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1614532237
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_220
timestamp 1614532237
transform 1 0 21344 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1614532237
transform -1 0 21712 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1614532237
transform 1 0 1380 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1614532237
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _56_
timestamp 1614532237
transform 1 0 1472 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_30_28
timestamp 1614532237
transform 1 0 3680 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_20
timestamp 1614532237
transform 1 0 2944 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_10
timestamp 1614532237
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1614532237
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_48
timestamp 1614532237
transform 1 0 5520 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_36
timestamp 1614532237
transform 1 0 4416 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_14
timestamp 1614532237
transform 1 0 5152 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_60
timestamp 1614532237
transform 1 0 6624 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_29
timestamp 1614532237
transform 1 0 6256 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_84
timestamp 1614532237
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_72
timestamp 1614532237
transform 1 0 7728 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1614532237
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1614532237
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1614532237
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1614532237
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1614532237
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1614532237
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1614532237
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1614532237
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1614532237
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1614532237
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1614532237
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1614532237
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_215
timestamp 1614532237
transform 1 0 20884 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1614532237
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1614532237
transform -1 0 21712 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_14
timestamp 1614532237
transform 1 0 2392 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_9
timestamp 1614532237
transform 1 0 1932 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1614532237
transform 1 0 1380 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_8
timestamp 1614532237
transform 1 0 2024 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1614532237
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_26
timestamp 1614532237
transform 1 0 3496 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_9
timestamp 1614532237
transform 1 0 3128 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_50
timestamp 1614532237
transform 1 0 5704 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_38
timestamp 1614532237
transform 1 0 4600 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_26
timestamp 1614532237
transform 1 0 5336 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_13
timestamp 1614532237
transform 1 0 4232 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1614532237
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_58
timestamp 1614532237
transform 1 0 6440 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1614532237
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1614532237
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1614532237
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1614532237
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1614532237
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_131
timestamp 1614532237
transform 1 0 13156 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1614532237
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_20
timestamp 1614532237
transform 1 0 12788 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1614532237
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_143
timestamp 1614532237
transform 1 0 14260 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_167
timestamp 1614532237
transform 1 0 16468 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_155
timestamp 1614532237
transform 1 0 15364 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1614532237
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1614532237
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1614532237
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1614532237
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1614532237
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_220
timestamp 1614532237
transform 1 0 21344 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1614532237
transform -1 0 21712 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_13
timestamp 1614532237
transform 1 0 2300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1614532237
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1614532237
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _27_
timestamp 1614532237
transform 1 0 1656 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_32_25
timestamp 1614532237
transform 1 0 3404 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_21
timestamp 1614532237
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1614532237
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_48
timestamp 1614532237
transform 1 0 5520 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_36
timestamp 1614532237
transform 1 0 4416 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_60
timestamp 1614532237
transform 1 0 6624 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_84
timestamp 1614532237
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_72
timestamp 1614532237
transform 1 0 7728 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1614532237
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1614532237
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_117
timestamp 1614532237
transform 1 0 11868 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1614532237
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_130
timestamp 1614532237
transform 1 0 13064 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _26_
timestamp 1614532237
transform 1 0 12420 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_32_150
timestamp 1614532237
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_142
timestamp 1614532237
transform 1 0 14168 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_27
timestamp 1614532237
transform 1 0 13800 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1614532237
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1614532237
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1614532237
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1614532237
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1614532237
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1614532237
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_215
timestamp 1614532237
transform 1 0 20884 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1614532237
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1614532237
transform -1 0 21712 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1614532237
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1614532237
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _55_
timestamp 1614532237
transform 1 0 1380 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _30_
timestamp 1614532237
transform 1 0 1380 0 -1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1614532237
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_17
timestamp 1614532237
transform 1 0 2668 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_31
timestamp 1614532237
transform 1 0 3956 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_19
timestamp 1614532237
transform 1 0 2852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_31
timestamp 1614532237
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_17
timestamp 1614532237
transform 1 0 3588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1614532237
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_47
timestamp 1614532237
transform 1 0 5428 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_36
timestamp 1614532237
transform 1 0 4416 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_43
timestamp 1614532237
transform 1 0 5060 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_25
timestamp 1614532237
transform 1 0 4692 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _51_
timestamp 1614532237
transform 1 0 5152 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_59
timestamp 1614532237
transform 1 0 6532 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1614532237
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_55
timestamp 1614532237
transform 1 0 6164 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1614532237
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_83
timestamp 1614532237
transform 1 0 8740 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_71
timestamp 1614532237
transform 1 0 7636 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1614532237
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1614532237
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1614532237
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1614532237
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1614532237
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1614532237
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_110
timestamp 1614532237
transform 1 0 11224 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_105
timestamp 1614532237
transform 1 0 10764 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1614532237
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_24
timestamp 1614532237
transform 1 0 10856 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_134
timestamp 1614532237
transform 1 0 13432 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1614532237
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _57_
timestamp 1614532237
transform 1 0 11960 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _31_
timestamp 1614532237
transform 1 0 12420 0 1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_34_146
timestamp 1614532237
transform 1 0 14536 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1614532237
transform 1 0 14812 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_137
timestamp 1614532237
transform 1 0 13708 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_12
timestamp 1614532237
transform 1 0 14444 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_158
timestamp 1614532237
transform 1 0 15640 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1614532237
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_161
timestamp 1614532237
transform 1 0 15916 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_16
timestamp 1614532237
transform 1 0 15272 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1614532237
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_182
timestamp 1614532237
transform 1 0 17848 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_170
timestamp 1614532237
transform 1 0 16744 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1614532237
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1614532237
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_173
timestamp 1614532237
transform 1 0 17020 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1614532237
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_194
timestamp 1614532237
transform 1 0 18952 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1614532237
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_215
timestamp 1614532237
transform 1 0 20884 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_206
timestamp 1614532237
transform 1 0 20056 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1614532237
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1614532237
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_220
timestamp 1614532237
transform 1 0 21344 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1614532237
transform -1 0 21712 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1614532237
transform -1 0 21712 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_11
timestamp 1614532237
transform 1 0 2116 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_3
timestamp 1614532237
transform 1 0 1380 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1614532237
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _54_
timestamp 1614532237
transform 1 0 2392 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_35_30
timestamp 1614532237
transform 1 0 3864 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_42
timestamp 1614532237
transform 1 0 4968 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_33
timestamp 1614532237
transform 1 0 4600 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1614532237
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_60
timestamp 1614532237
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_54
timestamp 1614532237
transform 1 0 6072 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1614532237
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1614532237
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1614532237
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1614532237
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_110
timestamp 1614532237
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1614532237
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _58_
timestamp 1614532237
transform 1 0 12420 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_35_151
timestamp 1614532237
transform 1 0 14996 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_139
timestamp 1614532237
transform 1 0 13892 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_163
timestamp 1614532237
transform 1 0 16100 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1614532237
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_175
timestamp 1614532237
transform 1 0 17204 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1614532237
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1614532237
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1614532237
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_220
timestamp 1614532237
transform 1 0 21344 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1614532237
transform -1 0 21712 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_14
timestamp 1614532237
transform 1 0 2392 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1614532237
transform 1 0 1932 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1614532237
transform 1 0 1380 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_28
timestamp 1614532237
transform 1 0 2024 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1614532237
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1614532237
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_30
timestamp 1614532237
transform 1 0 3864 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_26
timestamp 1614532237
transform 1 0 3496 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1614532237
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1614532237
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_63
timestamp 1614532237
transform 1 0 6900 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_56
timestamp 1614532237
transform 1 0 6256 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1614532237
transform 1 0 6808 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_75
timestamp 1614532237
transform 1 0 8004 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_94
timestamp 1614532237
transform 1 0 9752 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_87
timestamp 1614532237
transform 1 0 9108 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1614532237
transform 1 0 9660 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_106
timestamp 1614532237
transform 1 0 10856 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_131
timestamp 1614532237
transform 1 0 13156 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_125
timestamp 1614532237
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_118
timestamp 1614532237
transform 1 0 11960 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_7
timestamp 1614532237
transform 1 0 12788 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1614532237
transform 1 0 12512 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_143
timestamp 1614532237
transform 1 0 14260 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  psn_inst_psn_buff_30
timestamp 1614532237
transform 1 0 13892 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1614532237
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1614532237
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1614532237
transform 1 0 15364 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_180
timestamp 1614532237
transform 1 0 17664 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_199
timestamp 1614532237
transform 1 0 19412 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_187
timestamp 1614532237
transform 1 0 18308 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1614532237
transform 1 0 18216 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_218
timestamp 1614532237
transform 1 0 21160 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_211
timestamp 1614532237
transform 1 0 20516 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1614532237
transform 1 0 21068 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1614532237
transform -1 0 21712 0 -1 22304
box -38 -48 314 592
<< labels >>
rlabel metal2 s 2042 24202 2098 25002 4 ci
port 1 nsew
rlabel metal2 s 17866 0 17922 800 4 co
port 2 nsew
rlabel metal2 s 3330 0 3386 800 4 i0[0]
port 3 nsew
rlabel metal2 s 570 0 626 800 4 i0[1]
port 4 nsew
rlabel metal2 s 7746 24202 7802 25002 4 i0[2]
port 5 nsew
rlabel metal3 s 22058 7080 22858 7200 4 i0[3]
port 6 nsew
rlabel metal3 s 22058 15512 22858 15632 4 i0[4]
port 7 nsew
rlabel metal2 s 9218 0 9274 800 4 i0[5]
port 8 nsew
rlabel metal3 s 0 9256 800 9376 4 i0[6]
port 9 nsew
rlabel metal2 s 19338 24202 19394 25002 4 i0[7]
port 10 nsew
rlabel metal3 s 0 17688 800 17808 4 i1[0]
port 11 nsew
rlabel metal3 s 0 22040 800 22160 4 i1[1]
port 12 nsew
rlabel metal3 s 22058 19864 22858 19984 4 i1[2]
port 13 nsew
rlabel metal3 s 22058 11160 22858 11280 4 i1[3]
port 14 nsew
rlabel metal2 s 22098 24202 22154 25002 4 i1[4]
port 15 nsew
rlabel metal2 s 6274 0 6330 800 4 i1[5]
port 16 nsew
rlabel metal2 s 10690 24202 10746 25002 4 i1[6]
port 17 nsew
rlabel metal3 s 0 13608 800 13728 4 i1[7]
port 18 nsew
rlabel metal2 s 4802 24202 4858 25002 4 s[0]
port 19 nsew
rlabel metal3 s 0 4904 800 5024 4 s[1]
port 20 nsew
rlabel metal2 s 13450 24202 13506 25002 4 s[2]
port 21 nsew
rlabel metal3 s 22058 2728 22858 2848 4 s[3]
port 22 nsew
rlabel metal2 s 20626 0 20682 800 4 s[4]
port 23 nsew
rlabel metal2 s 16394 24202 16450 25002 4 s[5]
port 24 nsew
rlabel metal2 s 11978 0 12034 800 4 s[6]
port 25 nsew
rlabel metal2 s 14922 0 14978 800 4 s[7]
port 26 nsew
rlabel metal4 s 18117 2128 18437 22352 4 VPWR
port 27 nsew
rlabel metal4 s 11248 2128 11568 22352 4 VPWR
port 27 nsew
rlabel metal4 s 4379 2128 4699 22352 4 VPWR
port 27 nsew
rlabel metal5 s 1104 18741 21712 19061 4 VPWR
port 27 nsew
rlabel metal5 s 1104 12032 21712 12352 4 VPWR
port 27 nsew
rlabel metal5 s 1104 5323 21712 5643 4 VPWR
port 27 nsew
rlabel metal4 s 14683 2128 15003 22352 4 VGND
port 28 nsew
rlabel metal4 s 7813 2128 8133 22352 4 VGND
port 28 nsew
rlabel metal5 s 1104 15387 21712 15707 4 VGND
port 28 nsew
rlabel metal5 s 1104 8677 21712 8997 4 VGND
port 28 nsew
<< properties >>
string FIXED_BBOX 0 0 22858 25002
<< end >>
